`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
LzlnqZG83iTTWrIOOlvfzB6oWUzctHa8qGnVw0QwSLH0S5V+glKMpJKJ253ByiLdxeinZS/d+TXS
GN8wGYI5ow==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
sXgpoAbXllrOLkTkX8thb4wE/iIXrvnZtcG+aCHAa/Yc6J1dwW0z+oon8uvfGz6ZbLrzvrWPR67U
ONSPy1dhsM+4CAJNdMQIkYfdssKPla2TYJ5ArB42wJZyclNCkDyDJBE5LAxyke5BdPYFCGbq8V5L
0TQJe7pnZsaZWQfil/c=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
JuzuL0d/kwI9T6ioixhhhKflrXMOCAq742liJvdiTW6ac4+6lFkqIbexwXuEcPCmReMGjUloT2dD
HMLJWQmQn/3hfbDw3bawoELFJAn+leU0SgSXXOtjmwMq98wj9gSTPmWsl5M9ZMezcZVfk/2bRi5r
xpBzxJhE4MXTanmdIJOYxCREDRMADZ7WL/K95P52wIt0hisQSSH4jhwmz7/1u5Vwh/GxJhS9zGMH
Up8qj3IOaW9kJNqvvQ/ymKpyKOzEtGAQC0XsI4VhVVnCecA0gYFGocV9ITVmYW4ucMJDxS5YbvIs
sYl9mLn7V0QZKDqp+lxsCzSz96fPzqW5gweqWg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hGxCciHGNXd3ietLZjlGdou/vGxeQDo1KF+KIWwhf85ZA2+LPCRQTK6wGuFH6cxdDugQLG8mE09U
OoCfVvftIr8yPWi8kmxWL8nXpaXvTgsUQSrAdcVW1QbsB1rA+9bJPwRaVG+G/sRXStHdu9hcs3l6
8K9N04mDpMRVUk3w/P+xJvoBeQTIa9nrRb0nO7VAFoJZCuA4t/htU3Oh2/F9LMeElR52s355ir+d
TfWKQkCvSme21PQkLIrdm7J4NcIj6D65V316ACJCCMIiwlhwYTuHXAiK3nnYETQEqPIO+NFnAM/b
c0PhEnROFvrOZbgxbhfG9F8p8ZoTRpXo7oAX6g==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FmAbNjWez6M1NE2Fh7pg5kMQpPDHyB9aMNpIT8XyEkOHY7q3eFUAeFQ0lZAIGrvL7kmAIgIbodlt
Cmbih5loHgtj8M3B7AtqgSLcZE65DU3SpF5gGl8u0dJ/J/6Rf5KClqMvpAyCDqQcJ773A9Db7fxu
/CSVVEnKVrmbWuLcTSzpr+RSL8YyIaHk7yGVZuZyyZwoLXgZcu1yiBFygAw9p8rST40ijm+Z87gw
pTGXvunr0fl77J/vNyQwjbA/QJ/nsqp4TUe2KZhyRXNCchRus8B5Fmgs55M2byOMW+6v7+z0uFUT
LE9+EmbMtVyJUeIqSiJgvbmyLJrfTFaTdecW4w==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
nqmlpCLnFrwo+JtMnJfBhSlGE2In2Y7hsJp/sqhZ1GkW5+pyc8MDjSL2mfvouEbSWoK2JH0f71Tk
tPzMEHwz1MjLYiQhc1YrYPGbq2qBm3ok9dCQXGFZCVW2Uvo+FcGRAns6vMHssJ7x4HW4bRsvzKpw
83lC/s+ZTdqign9s2wk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pWGEBayaNrx2z/G5sHCfeu6VmSrKVbH6RQXf/i4Y3tQO6hCI/KsXfho4nsQKwhCB3xiZXgXtnSsf
sPATlQszo6cbr5TmIa9S3vs/cdztrnDNEctId1iYNGNxedRd6+7erKh6xN8bU6NY60VOlm1BA1bS
wC393TAerqmp3UIko/LPXBdpPkfmomJb7vEO08b78aDryoNSbeEOepayzFcMzbHS2fH1MNoFYnz9
rv/FVe8O8j2YDlv5P4HbrdUhdO55lR6aI8mLFX8A86sAqHXzcdvuWBxpLDkbUBFxV8CQoKPvBIUl
fePxraqADXTB1CR6heJt8tJ9lTYNcdqX9NjClg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 246912)
`protect data_block
Vl5F44U2/61F1UUMTngMkCpgYWHwnGMHU+pIvXM2kaZ05Tydu2wzI4hs8mL6gSwOFksVfVzIPfan
RmTNXe+XJZU16ZBh6JfexD9gf7srzTaWrInnxVramYvlsrZs8pIB25M8khsF98KZ117Q0JJnl//A
vF9JfzIsLC/i+2x4m749qZfIrTSjjtlUm4iOop0CnKZU+FlT/Ra2Ly2aZbTbhchjQ/V6YQGiVfIr
m/dqeZ6aEzzOlr1Rpn2fWWcfFaziWGCeF3TTog+zjUNQYWmeVJxFLx65ElWwOKB1rbn85VH3Wxcc
XDfUJ5su0xJp0ANoT9Cc8Bjm9NM+RJXRvLh6H1HguesJ6nPG7LiBIuZNSE2rPbBinX4fydZCmk/C
o3hZoOs0cmWHA+z2XcZS2ahNGMUrsXEm0sgEqd3b9S/EDIIA4zaZbxh4EL806ojomYnVj5VmFHUq
dWr70ttNuFyKs0aSsKY0P7puEb8glPkwYiGTgwhwvvuDjSmqLo6myHF1EsE+xSmApGmF63dJWFv5
f9/HyfEXfIcos+pKcxudMRcZENos6BK7YkyMsNLNZgEWlfsHXWe2fLpry95utaNc955RAdy3mfa8
La/XhmKDw4mKiMJ3toTcOgTGsvd5W92IaAWhcBurTl2lXNResvrYCjD5aBAnjFqxB6jW+3LAX+5g
3pbDYGgOEFbRWrykOItkxvNhJdvcRnO/F8F+Vwg3RMcMAn0V9lz/fXc70mVvM5S22CbiVK5W4duB
XbuglMcqN/TsRPhhZE+yylWRR/1jNEjUV1ZYjBOjIVhNgo2SFYfNV7aqTKnTM7UBknEEVenChPyt
iHfeY0AcGc2+4xlAIh8RjLB9bqOjkPFeFWmXCJhyFSrI02yn7UzBFhzuModdIS6VQniM49IqnVv6
Vc1pRoBs49Te0sFgde++HlHWvRl8VsAatVBSTZiXzgulRc/Xb5/BXFpvx6BjYE50rdCzQt/6HpxT
zsZosPAmbIaCRYoEn36tTBeTxQ6cFRmy74/8MKRt/eV4nB/OhMEXeepnltXNWUvjLjPivZNxyAx9
uulSxDEkCxVAY4G8wnv+PaI2fTVgZHuhbVnpGSh1B+7e9ZigS7Hx+KbLqS4l5L/vv8uSvSMORHEo
rYjEZERAJV5nUauFKQZVRShqe3zoc1tdJWsSSlxTmVNBp1jGvt6QRvFO0wgipwabBCwGHvZXdHpg
yY02JZa52QaGnSFtQ7/e81gFxsmTNPctZQDuQJQ/XveYr8zlbyTmr075nPNPp4sjFzfklyLGLQXn
iSoT9RGjfC/57P7A7H9sl9gFs3vGe11nmrIHLQRLoW8y7ZlZ7HXCjGyZqNQFQwawEpkvjxmiRa0r
OVlQ+urM20353+pPHyq65NVtVgRhw5bm/ZEusVjJTinMMKey3K0U2JTLzNhdNvD11GCPOEk8vmgf
iJ3kFlWbbZTreRRrVVZOlM2pXCDDeu4niuWuDDSXgI9FLERoH31m9tPcik2zYjYlpbC1+94SO1GJ
t9jCpa9kw/l6SPwHapKIffIjYZQN5H2fnCHKdss4flGA3bmE95hjf+v7l2LcKBctPn7zBuRlK4vz
D/UIJU/IP5uuD1uL8gXgrRW09Vjkx1k/iVuC9Q/AhwkY9bKByOosAiklxrKZU16rEbrMFMiEDvXp
1WGgMX8fzm9FfstngmeZ3QX1s8tOk6aWoIheDBkjd7AOqfd+S1xjGCH/lrAvp5wEcVBfLvSH+PLn
AGdgSdsNLm9EZgkuZ70MN1xqkE7O9iX3pP118P+2GmORptOIHlfDuv2XyNcDQa3jeFrOpi+Kcfb4
0sBcC7rC2/XJbuJnuCdIi90njIEyRLGXGIjSMrhb0EUxIst17HNx13IXkixi8jiBuTD9jiZ1Ud1g
WaYrbbkLfUf3bP7OUVNE8Zl/HhQpptgHiYinQ5CFkxnPns7CK4zbx0Q1YiaGiKAtXJPe+uBbOkoU
+S4BL3G2VY5q+Juil3Ge4+GwlqAQQk5Jaj6XnULEspWkLcCBPfgHklExNlFUb+MvYjRpm+mEeBHW
MrjZUoOcQgYu6JT1repaO0NOuIWb7fxDZXwjCOth37W3ToO0C3RtNbMaOFpMjqIJBP/f2ZnghdE3
znSZX+jqKOOWGPcNQL9fSCiTIrig0fxZTQn4pp7ky01lIlqu5TTwPz4PY3CxerwqA7P327nIF98m
5JUx6cIiNI+3SuUkYbhfCPHW81Qja7QCOQeNPSsgub15c1kDH0QwUSUbkOY+hovoFKTkI9IXpt4z
AiqNPO2lhk3i1yx3OZGEt+1n6x5CiRm68Y97/nHRINo8YfRRnXGviadDmxFf1NLSwghXIp9ToWWX
XrnqWLoiB5TVjzmaV7smbrecckkCPSFVA+NuR7K5PU1MZRn15eVCv9pMAPqC1765l6R7hDKdFxRk
jvGbwXF9DjNCfQU/tvyLcRfuMCJNs3BbktgQmonSfh5sVYWbsXH3y+kJIJonWbVo1FDGLZpnrQNz
2si5w6qmyetr2kpxxa20p/gmXcGg4yugfZ4FmQk9d4zPNhGmpPgnQhZkciYbxsX3cj57m1iuTxu8
/zCgMgJbwdGzAvee8kS+owL3ZNRbKJRVoFhdB1pZYKCVxbaoR2OIKkqpq6V5/F5QfEfOoEpRXKU6
xDwOr4gnk+wVdz6/VdCYfI1M1xn9uz23KXoDMU3vL9ucc1inPX0TjQXqz/zEq55/DpSZipTiQlhY
gxWQP/DPfp+igYdRC6snHcgHDEYNB5MbBkYalMYT7nQ+9CqhL8UJajpxkklLT41rkrMVSwbQZJjh
BtJNGlY6SnbFM/T9Vjp9yrnmMqL6QPzczlsCWu9cbDJ9kpKYB5+LvRL9JxyT3XQ44+1wcOmJ928x
Ye6IgJb907RGnJFKRSgxILLr/myGmDNki0+l4IlQA05AibaGu33m8VQV5y2MaEo0Zy3xbD3TUnQQ
+gimMlRC7TciBM2QLedZxC5EreUmRi3g6BEmbWPKsgX0rrV0FBCr0sVURipRBphS5HM8kEWfYHdB
1W/CPv7AejtdTEqoTMm+EGXJ7vCbggxOQSsLMoSopkc2pSzgTWdCD20Q22w4AJSFkj7GYZCqYH2J
L5n8UfjFygW0EVALC6M39Et7Pgxpr2q1z71dAc1FY8Jx17Qbc3lApVFfCFOJxXtn/i8cttYNXSuU
7ZRobCXHMAhw73/Av+XDKgK5mzKEzdhif6RdID78rIi9ZB2zkDjYHcITeddS+Bo42MwB4SjufBqE
KpfJ7dKdF8qJyfIpmEvT41GMuOrEn2Ls/Mi6KKpzZe0pbc8CmSxxX8WekCBs3CQzDGaPr/riMZKW
Uz6lTO6uol2MNHeqESleqtfavXtOKvWauxJMc9BwWulq6mJikyq0uLUgrcrXAbARbQJFLwC2A7zh
roIxwTtP8rR2FPMkI1HEwBwjkdNFzrcjpqnG3U39c10dxhLb4M+2DbHEG8aAQlGZDPZYKCmwTUGd
gRqiV4hsg0m7gdy7WoLgfPxXqvo0VcBzgPXj4EU21800uj30dxXkuMEa71A0EbKOfCH54cEkiTS1
ajj4zwIaQgAbMWdihv7CCZyNdQrn9aEqhoqj5ai2OJuv1wrm4D5Mrg9AOW1J1pW8Wy1831mGzrGk
gNKESsBfV5FtOEQyjVRoS3q9Z/HBbVP5r/SrWdDQ3e0ye7f1yXrDJXHxo71Xgx8F0OxKAB4mP+OA
uzD3sVLB2cvQm0Q/o7OeZpWJv/f51b3OnHrRA+aRC+/tamPyPmUgxAkwLfpUVK8caKyUQkhiYB1e
XZl5dxLbxsfhALokwueSCtJHL7id7dAx6RhaVrjfTRtx6R0JrNID2/MFDM9dcV8tdqvXuHvJvIty
B0Q07AHCKGe3CezwPtMi0STggKpyDwbMjlocykmOLnn5gJHG+nJIWFmxTRJgST5CD5ytKz3BIk3B
/sI4CHHTFiaAKGmwjf/x9mycslRlvmP5xkRH+3CCEC4JEkNhg0Dw7v+skbWXomw15lfGS6eOkOxg
H9YutF1UtLu8cv2aPPirjL2IXE2m9noOVFl52PJsXMZ9DN5/VGiM6KcIGDnxwDtxFQs90dz+iZsT
SgFhKmAruRjPo3nIPWGMM3Jb6Lpl/uG7/Mh+wRPIaH2jdQj7NBfa0LzJfw60QG66t4LZBhmUP3Fy
IBCp7pNn9gqF15MmFKF7HUAmhF4Objd24U5GGfwPBep6lrVtCHNuOdL9BZFNFDtFPSCSinZqHYtL
jUn6ZyO3bmqVIqy5cHsyuY2Epzj8ol1IhH8So29wVWxK9EkiOyHth36ohBrfSletJyMjVdtdMiMo
N8j4LeaydcLUAs9pCV3rRjSWVFgImgvypQlffc+J2KUI7U/99pt1UGFsfw4dgC4h/JMlKfydAWmp
tjTzzZEaK7jWXEkj31sZqHwA1IoGEGMrBmNoZlJ0T3NmkuHv4n9OJdmIwuWyC700QSmJTrrEYfug
+kdkNrYQsjmok3gRzhJmIqF9E834trgjc6U4FP4kBLartcRwmqj9PHFEnOYHZm2HkblHttJOlm0Y
W/NUlV6NjzadSwQibUqd4kdGgZBd3W9StnkwyofGx1WRuOf6Kwf4GW8zQCgKPU9PjHTvw8bi8ngt
QZWatoT1drUrwKup+aGyUAcWSZYUGs833j3HvoXWXhjk9rMIdIapQG7PdF9Y5ctzGGcOGsJuveoa
HjspI/MKM0I2ZXsUxQnlTOs5/GaLpZZCdv0uYsmHf83wSDyAXvtzcBZ4r6XPVf/bH24IMeqV03rh
w5AEv0ZF9rhDHnbDqj9yCyTElvdQoCPo1tAZHWcp596LscfeTx/ZG/SR72p/lWPOKDlKR2gL6T07
aOeJkpPwmq1zxjGFsfko2ivEyLCd44tWMfk7oSgGsno/2+0dSjZyRHQqb+AplKcqxH3WhI01UBfs
GxCOnByYkJYgMIk9YLZXWIh4AniBljPLP7DpHhZmAXp8CmgVA3DXi7SrrYpsbBpAf7AMpN/RXKEh
McNJxzAkvH8iOsUpWr2F4vcUa+1Uf8AVltMCRpEgD7vtFwwh+g6joc25DLebf3oHJ12/8A2/qEZE
GHlSDX2Uh0VGLO2g9g4rRVfJd22McDJXg0omdVhf2tET7xlDVr/QulazKTlV4DFLcwfI2bVyS8//
OeFXE+EU5SqYlijyVhXEVHheAzJqut0zC3rkNK24OTKBqt+eXyyV87TEVHK+ERaX9dvNn4A9yhx8
2VMsua9zOrrn7JbGdYnNX0Wp7+F4rNh/TpLxGsEuaCqJN6B5c6D3QPxYzg2ehJWFOFFduzjXD6jQ
SCHEGxBIX2XB72s3/ZQL8KsDjadENNLqaQOP0P7Miy37Rk5kF8MnBlY5gzgrh1w1xtwHKCJTX2t1
btXfvLxdne2sGQ9ir6884qMY3WOLKys9kayodOfsO4a5hySFFtAxrilOf4VJbZTSKfejchKxXAse
shPL5Lcebmf8Vd3tKdWorjMtppaeap2yJCJPOOReW63vaRAX7X5eVosABxTUiE2ff3ww/PRF+qc+
CeL8Jc0hxybZ0fF3eq2stxGXJHnyHttCnQTXP2mXtJ8GSYOyhaIIb5li5MNtDbZiOsLH5Ed16o/m
s5Hsg72fFaZgt/o54BwNE8GXkQGWd4BeTyivuG9vY9sfbqrYId8vPJURarZRW8eaAnaVlcJuvtfD
AP6EZXVz5cEgwMX/3GQkN2ysOOhpXigZTOmgvzI9MzooB9QMkeM2i5NZlboKoSkm+UwgUo0mrUqY
NnfnI2Qfs1TRrqtwaTaaa6yvrhBBFtuZD4rU7ToTopBPVzFvz+vEUXLwvfA3fDe2K8LuJUxiWTc7
se8jsBIePCZE5UBlVSnpaCuZ5OLnLDv7uchAoCtknvB4JVvNXRqCaW+F/FHpQmeasNA7MZg54ibP
yn3oG2AypJRs2MWg2nSbvb8JUFBjXfh0L/nz1VlhYL8Tte9TLfZKzEWKLkOQlA6ohfnkrNye2vl5
2CriZOiHBo5s00J/i5+teZAzZb1MZm1RQ0sbTfkqrf1hGrUOhNoHaLyXZca9hWVxLf0ZGHruaHfe
4SYDmrj+VA2Y2us1Z/70q/RHezCTAwbaJz4HkSSt4C077Kjc20kO7Ts3ZU57yWJekUotdvlBPFpc
TBZ5z73QEAX574x2T+pZ1Ul9v9UQdBHfwbXvIcpJUaLRIxQe8huugRFbfUICKAWatZEutYtmCcRS
lR90RJWwqov4+cRFQlUaSpC7nsFY5owgZ3Yx8x/Mx1TCcoghTgRqsNh8OLhZmLiJddZy01d9RJCO
2z4jNjZnKb/eVCxloJ8nTzTMos0weps9Pt60GN4NUNk39mCpWmHLmVkBr8upLYhbW3W6K8HwWSYq
ALfTidEe4UStqX0BGaEVPfLAXlTtUVXpG2f3wHg4iIrfpdMK24pwhwZ8OCF43WsGoDNhsDYqHDiT
/06gvHN5viN/Zj+/1D+S31XPxzEnrO/tNNmOSyEYdUdkEmSv6d2CzwCAyr2uBtot5TSVh/UdwVUi
xRYAshJm+EXgsvriM71u9YhXwausPRq2Gq/RcwyyQ2gzTjKxlTE8/9ZiW1i+zvnrYMZ74XAKzS/8
i7LfjasYFEIpAUin+I700NMTz8FPSFmID4uIwvtLovLaSkvl0zy1ZNvNT3UQRLickD3NjAzEcDvW
Hl2+qVZL8JN6H4KV3ZkbSWeu+6OS5lIVnCMeWuGThjNSnoAWG3Ih3ptQmozzV9jvLalR83vMH4y/
p/mxCYv7SPCZZ3MUeO/b9RkDc6ySeX0ES4vfITXq5DWqseKn+FfekNgAfHYMK6S8YqxxE5qyPU4v
GiosbLFqpY+J+7ajjqfrCLzTfRJ0NomSqyU9AcW1wMIgRKyhRNmyMq3+lSTFuEz6+e0uoU6qfcKs
Z8D/4mEvJ08BsC/4I2AcpiMqOUepuwX/IHcHtIFp5rvDhSv9NXkTiV9p6AJlJr47pJQeIupawtXC
CqEf78u/lZraxUOPtAKeMiTS5Qtpmnozpf/glJgVqKjFDbKe8gCA6R07BmnjIB9tNbhCpAbdcj8j
j7DZ6wyW7UVnQ+r46dfWJtahY1ZeqQUrTwRToiFBsF+QzueGn+3HEzfj5Xv56N5kZ3OwbzdGJHoZ
JD4bp6xTgL/cyZa1Czq5rEn6OUDF3uDuTFxs5949WQzFayYx1vqYktZBMmJL22OyAtShG5LxIejF
+EHoApp2HC8bzubPotvHlgPj4BKn35/Q8x0G6ZnWteZY7fB/gSvKiFN8MQIGc8MK1yfob3TbzMNk
2yZ7625mNzIAOVTd9DuQgU82aTPrVeh/H+X9lS1f9P2WJ1qTocxqt9j5lApbE2wSM0OIb8IP8ENQ
Ta2PSb8Y5YmtLKZrzYVwdthpiwXt6IR3P6mJ9aqqoMrVpzfox8K1vGOlDbIercfXdrt9O5VyVH1o
VzuWCYHossadJNuXz7XkVgIIj33wQC0DUU9B6VEo+khdRFMn61J0mWm3geVz4Jr/o9C6V4Kx8cNg
FFxHpSR6AhPLl+28VqwJ7KAb2AoPAdbC/kUaXhD1GYxqASFLq/5ObuPPPkSHZIyTMVHDxkYyCkHF
Wtu5uchYSYvaqzLfO9BJn2H+7RoSHcW1AhPZQ5OjoU4YtTB1yUX4aWhleOskjdlbESyh7TCscCEJ
trb3rypHCIxNr9bjLb9hhIWAWxeNXjVxtjR8UP9cnuzeTd82cbLjF0+dD7W3S0aKcHqoHYB+HDEZ
NS8RxisXFz3MUAAW42uIshpXSgFsdXTpreq5R8TCRknmOFjOVzIiOahkscMpIvFVWzJxcZlItf/Z
VAo468fxT416gAGTDTlG9E+4LsOAcOzEoF2hXNn3i6Ps8bVNU7cg/OZkWp5cQfu6iTHxWztfXGs8
+eDZr7z4KNk0uqMUTBjQ4FSALDsCewEgNTX+qoCesTOt8FtXUcZgtKL2jlDWx1jJaGk56SDcSvwz
SQM2G6ezyOpbGV4j+klJNhVI/dScggWZuFsJJKei6G2JLpVp4jkCq21fjmH8V2BmaQqeFgz9zkTT
0Ib3Ewm2DITg8kZViiHJYEWQMoEkbGvlIwXb+NJDFOSrNoiG4+Nc/r9JJ4hdlxGfd5ybgEgjFJPa
IwcVWU6SZhioZoYS8cIhZv3DEVFJAHoDAjmQkDD8nQHaWXsa2r/ZDeRyn7npsRtIs2VADQFbkWNY
K3DQP5jZCl4+QvAJxNzem7Nj/jHk665ddHKNFYLOn62ZsPyxMCGC6jnxLgH3nRf51UEORHd6dHDC
P0DKSkQePTgBq8ai+hK3ekfF15BtCnT/Hlkl1qZ51TuosnXCC7pMWlruG3k4Y/xq7wRbkYpcQtPZ
vIeN55gifDheqzMQmh40at0G1wd9blHl8yh3Nlwb7HVgj7ESlTzepKbgx3PGLC8KXgm2AITsZtnX
pzNMdqjfzDS4LLdzm9WgF4MgeUnkpSWbS3dNvX2SSLeZJK21SNJ1xON++RTQrsdQq229l7cmijRE
13rH2QqrbL3n3TnTGFswg0fKdfCF5FNjo2Gl2XrmpOh3R/hwNJLt/1wulDEBFqdEWtHaHF3oj9cp
W76/mpBtUwp4PoPPRD5gLHcf7pxSM5ibof4ovse3/ajrRZGdTNrIs74nOjwVLMbZDIUKu2ZH/zip
Sh3xyceHu5y8WDpt5pKO9CADmDA1QdoxZRO7DROD0aryn2+h7WkS4eMYkgesqWlJslF4DAvO1ygT
bSqMHBxFyHdjOlXw7AUOsFeyMu8MfNTHxY45wzv1qvdpvEH9fruj6RxdgItpMn4OiTFsiJH1+eZR
3yGUhSZlAKo3XDcreau07rYMt99iSK6ddqOUqyhuZf477tpLkn9OvXu9FDhGC8qOJSb5Do9PmtxG
9Uw+rSiqmtn6sCTLFPF4jmM+SiT1YXlTpu16PbupIpWz/WHx+VCaSXJeidffZKYeFEs+WMuYUal+
x+NEisxKWcgep/CSEaNHYAOcz8hF7rn4ubail1664v8P52QJ6D54RggV9mIONpkzGu3RUkAISK5o
P6FDK6ZanYltkFnhpVKACAxhPJ2JWU8xI/A6P+4qB4ngzSbg52xL6HP6pGER/HI2SCw4vUJw60a7
jMPXx68hAz2McswsD42Rpj4+7RGQfGpDe9Vq18bL9ZD+1gPramb4+zD1AXozm6roVwb27+l/ElW5
xpBVVc+AbERcK3Nigd2jKXfateTNpQDK1MV1z3Ebb5fdFztlWAnu8tFvbltSXJkziOYna+0JfTpF
UUufNyXsDrAkmpWzWSacSvIZO/X8Uk4sVyiBOOgQfNlPnX8VeVaQ06Wub1Z2eqkwTdUTxKzffBJ2
G1gZzw/ZjKu0HqcNx9Rkucj7mhrvJlfR9ATYDoCRLXhP3jZH9zrVw/ipvIIU2T95W7D1tWM/rLwt
F3Y60Aj94nXhSWTsB86TWghWbTMyBofCdqJJTsOBkiORX7Oqq4EIMgb4S4+JEvnLL9idAWgO/Yy0
MGNNtjUoEBZqZoq7MxOr36gYuogt5sQUaNe0LdEHv5Ij+ejEWYR5Vve4V6+ZoIZWkNtwcFvtWqzJ
J2vK6jrrQc4DhAj8zyd2YwQb4r3OaFNk23he4ur4nDXMlx9JOv5xrTehK+Z3Vt/7lDKv2hczV6VP
ZQAJ21I2EUR5suHwsq8VECdruNhTv9brynIr/fgKkna0M5uUGNgTQIy3wZK5PyqRuO9GIifOkv6d
vgZQvAmUUFzBeG8RaTyrlMKsbJ/PaCTKHsrmSYtvklctqFh5u4nomIreibH7AdW/rYd7JNd8pf9e
yvhPCXKIjSCB3WL5JZnW3Yu55QJLX4y3ZxQf8/HR9W1X5bEcKZNnLalSnEGV5/1HVjOPcNdpI4SG
xKnp1YTm4+PiOW0ORmph8rHql3EGqNM5aPeOXuEXjpgN6EzZ8KeKW7Obs0aCGpwupbVu5DH7Di5h
4EZ+6444trqsnjHLLBO11dtA9xPO/Hiq1hp876/K2574777e0oNr3CNRFExZE1c1ksqcLQOZJqWg
II19C0aNJJwzoHIlCTrRYmfEO0NYKEHAWu2WW8GN5cpD4nzYxrHKpe35dg15jpuL848NrtCBS028
uH9YQaxOtg1tfomzPs2uD8hQrA7V0uLaZuGTpZ+5m+BA40YmB3nCY63IbeG8WkLUZBwpeIIl+oO/
aehGZaAqnBiQwO+e1KMUWaijdLKiHqIKJh5lX3+Q92DmLu0BR9Fyeu9lx7YdRzU6+7s+UhwindCo
N+nLfdgTNoWt1K+DWYg8Y5uh7cRnEUXwsNG8yEivs0sOJzDDi9N1BLOEBJXzNdQpGfBhdFOrobu4
HKGBc3z1ScXJI8UdLjvAmxTmKLtcaqFJzZWzEniST29r8ijJYZeEApyRSN0C9GzyQP+wSPjDShts
OLLJBParpxEtjYLtlA8hAHLrOTHG54xrF7lqUSReU0bQyuO7H4i/xxbI6+ivtjKJbXCZB23ETSFv
4f4deDRpb0Uioonu6vK7cic03WdOjCX4QbEcc1+ojP9YDp4BeEmhqWZ5AdH+ytWxAIl/o6i+Adlt
iAr8eoX+aE/UytjaCx6mbPPTycXbuzw+awXb4l1pOF/mbjddHRaJgzGIm17Ru7nMQBjOm5Uyqmrr
BU5dFGDTmHou4lR3f2ipbzuQw5Xibtvj/FUa5Xqteg+fr4XboJD2EX/FUrvGBUUqRxNdRQA4z2q6
HiRxPZrtczEK3nI0P5WfZD1ROz8R2DzoqpYYB4ZjOG/Tks4TWdSHyH/9T7BviE6EN/M8M1N21s2E
VCqAKBR+J+dhTh0J1LfWmbt4nHu+gXY9V4RC7vzCfMKFjAZ1DWibSzbPl4MMG7mL+h6/DOQeBFpx
ijJv9iPHFRjT1tR8yzsYrhH+i7poGr7HcD9kqHF5u2S+YiRHeQsxGOS569f1HChdMZU11mO9i/4E
u0iawv/aJUM2rYEIPPKSVgmrfovpt8tfj+HLU9yeOzQwyhv/NbLmg1Yuo04CYwQbVV4JLDH/HuFU
v4n8WKQLL/ViuulA95vki+9WPKMnm6K6qWEoTVCBTcAf6EfXISvcl4FLKL7Wy77eu0hFrMFpvkkx
9JTwi2PZBknSoMyjeYyaUABJQU0YWtom6WKAB/dUZrKfzkQkbvDP1+lAObOY3XCtuegg7t5vhu+U
m77bzRvTRUyTeTDADLgBBJkkjvG+VxQWRbxf6XOKlwLUy8jr7m8QU9SBIbb/m0Kdd6xMs5TkRWUn
31tN5xNrcUvvVGXNbZP0lpMDknOtGqSTOHB/5dd6hvSzk7FKQ92UvVyGL+tMLUOHX4b6g/rnK9tx
O09VYTuPhkt5wyh1g6cODdGZXhDLX+EeEmpH/vGn1MngsPJgHr5rbpgLokuNzxlN6H5GCsbcNNt5
ydypdDO5B/J0Moe2O41dm2FyUHe2ls/i49gDwQqe6MhAiNTIV88kPSYiakCxdTfJ6hc048Cu8U3E
WWNHgRUEIgsUtwknsP62zDdIE4eT772ybQqFceHfbdbBncCi21fUX8wxezluR2HYLSkPC03dOpyi
V6Bq4Z+4azkVaVTEcomUQoK8FJdtiDRUBWt9fGyru07Ipivw4BSR8gG0LJG+Utb0dnD71sbvIpPk
RHnioOkKQJ4NTWb/q+Yf3/iQBWVraQFMfV5oxpxm/oyXczN/zuNpo1rlNTNpHXazBxDCB2aHOGuh
5/L6SwJxgMwHgIdPKDjxAdLLJRHF5uge6yWRLhW0OOX6oBLzWH+j7Zic+nB3hzw5BfNUlvUWTMb6
ItGTlyv1uA/Vw3jmqSWayyA65r2WxNQ+OGVhC31WeAKfJX7/99z+R2CK8Ts62did9h/rZIXkJhDS
ODWvGcoNMMrkO7V15acDAc7A+TQNhA13aBoDI6LA38eeY6AQBDUuzVSC1KdXVKeWi39CZX/7n8gj
eVlZrRHd4uVK4c0kcyWnJ4cKdq4u3R+3JCVPDOYkFyLkoFHI4RNq56qt8g3lxtc07MiSZ5UV6ZEL
k1VHNn/BFsNi8Gg3dHdUt3KnubMsxjRS+QfwdzjhFWXZbxrWjvg+3dUjN8xrEKQuTPLzU7S12tHV
Vwt/OHSai+vNnKu0esP7R+/BmVBh0NTXbZ+Nmt59B7kddo0StoMIU0BIxJrFT9c68VdAiBYuB+Ge
YJ66lv2Lhe5nTll8ri6j2tQTopnNVtW4r6ar4VIBkuyBfmQs+AsBJKvHHklFnwxxxCkFBssm6233
GhErDn2VUDrSscHZDFNEJZ70Ekzb3z5xEvdoHud4nZfHpogb0JXgPTWHaFBTFC0/GG6gM5TIZWpY
IKilAINhpZDRRDfAoK+kDlMY9kh9fWT8TRceioV0TIYhSXrYRLXGkaBceY2PWMBd6jANPXjdHf/B
LdsVU8+r9UBgrX12zf+FdfCo4/+iha14316YJK2md3/ZIdZvWuGYnoSik74gV5jRT6apo7P0XIv7
dl2sbVi95SpnG6tDmlsEokHVEsYYYMK0y2sNyQ6eJ0LOryTgC3lhZoc40WNo/BtyzLtFzU4VvRh8
mPQkKUXbsjKzpm2b5fCP8gMDszRmsU2Nb0CZ+XV6KgPcI06LNP5pV1QdVH/QZTfv3zuRKLc7rAJY
NVIJbr4hGHgbmKKPm23iUJ9Df+I5OJy1l1GchztH5JZvRIQbhdqwmYxXu7o+4ecTnCurr2yApe5s
GkTTJMDcr9pLUqtQltwNCar04B2BGurjqkC4fjGnf2QezkTHFsrD2wNLJuzORwRLnIP76SwYJw40
BvprJN4pKfEBWeDWgHCOh5FrxBYQfalnYXHyyAXjcDB8dmLKhrdspWbYUc9RSWFt19C1PZgsH5zY
QX0dtynR8OHh7lZw6cpn516jiyRNXvPUZvgSR91CkXKF2VQy8njwcgDAwWeMqZHc5QXWpFyRSzXu
6GAxhYnuSsS7BZ7PHrIHfD6br3Pd0+G0g0S6Yw8K7HB4d/VxsR/Gg4x+xGj2QsdeZNwgDMCwYZ3S
2LrrSmFEuBIclOeX4FbmwkEbBVK4RPzVgb8atIKzhaNK1Fu9sTfwc48K1HjROgqNflcYQJcNSJ0Q
IFTYvZD1/AhSH16J7PgRi697uBgxsH10U3KWx4HFjcocPk55u3H7TGWP6+TOwP+Hv4QDFLc1oASI
9gakZmkeVqv90diKWTkyYH3RITbjgaayPMs49WfRMXdMZdtknrau99mbx+fPCmSq8bcAuW6ePswS
fjBMFH45V9xcbf3wstvEmQ19Wu3ODq1uWSYyi55g94XgqXpcDD93n0iiAXO9DjQkQlN4ywBKs3WF
XwhoO2rPTPRk5Ld+PEFyJiU/oHSTteX5uq28Q1UAWb0xVi178uUHHeKAkWcFd42uebX/ROuQBwKu
RtrXoL2+94s96+8jP1BMB1T4TSWPH+ZW31ysjgLGZnP84THgk/s3ZO+45bAKw27bKL9kqcdHH1Wk
TxL5PJySYtNchBtborxklDgFsQlLFh4Dfcn2fiwP9EmZSQDZmC0+UuveUvaWMyt4PJnCLhfi6iGL
eMdBe1L5p5mxgw4eUxr561AFcU7qD6JvQPoLtR9aQQP9VvT0SsVN76zWHtlzjHhMaihk6Tm3TuuD
zB00QyhjhllZZSBHOiB+lFBC78zH3qZd+m6YU1XhlEO19u8nSb42BZcfesRLR8MtL+O8ef2D0Nq7
h3AaR4YF3zEoGSE/sn6IB5al5h8WIP4ERKy1XJAB4V/cLJFhoG+Ldx4RR6b9J69S7wd27ijdlSDt
3aJd3wYU6/SbXsUexgetAThPHkJHnlOHaXt40O5lfhMQlChpb5Oo2GPBaf1qeJEodxLO1YscrkF2
fIqmBfe7woezkSQXCUYp3Ghdpn+OnAGLa+5PwaKSq+PT/OljBCujiuDcHKC+Qemc+okRr8nWwf5h
Lii5GHOaqgIxkukeiDr2Iy6Zv2/v2VjznQqFhHbZA1y0DLaJGMhZJv4wgo/JEkVsFyb6f5dIdAfk
/mBwKy2sR8W9M7efTjcbCQDpFs3wvcfJd6ofJ0p3PJwFFUG48ZqN7DPic3TN3pUkgr366+i8Q4GZ
aZxYrTlsnwaliBZyjjYiJlqUbMCmRYM9lldvf8rCn58ddxWG/BFdHDxWaw0tYq+nHf9XQaGxpG9U
0M+tnMvA0zvLn/1lUHJeOkMHTgwZeEeUmtKdBUYgUsgpSpwPjYU3GbE4Sj5MRbOK1AlFCVFhz/IC
2kc3/WBOP/Hpeh76QmC25bU98FU5eqPuCXynJa7883ttJDwW+QqgrgVfDBTuw10CcFoC56Z2LIN3
XuLlNrH1Nispk1ZcYadJB7k9JRZ5TUNJmnQ4VwMSlsC88Ikeg6T9RBcQ2bLcdR/fI1N7NgoitKjn
l0Dn3FozE1pbadtCmjiTUEiX0NwV00nQ1hY+LuqA/JmazEXoV3UIgJYMqNG29INPJs/4DwvsU9Ft
7/uId5e38trm5xiyjY4rjJtUWmIHrrQVryL5JvynFO4oCgQgADRSyIIFx0iESyEZeWAAxEr/rm4A
tFDM2BBhry7I6MF+ZP2pb73HaTZOp1Bua5VKag6fdNMawJCc0B5GAlLvzug818E/+okbwP/VnRAp
5H2jwJgjdCwCmjGIDRDaWwfxJbaqfeM4imVPKShMgJ2mnyudx4DzJzgZcPZXNdrSeN7nICkYRygO
Nu9gOJGRZ3npJzBwvHCyHzQLBFAaNNCNaNziPL34jaKw/e89B/L1+1bXbBySRjoxC8q3R+RjLC5i
xjGS+MngoRT9zJOpoYp9U+dgIkpWqZYOYdZA3nucewOjb7TZkryG+5JyQAkawr7cOp7t0xNBrOyL
cGiAxIo78WU3OCOnb5WYaUyyGpOnx2b8ELJzsS2nkkXDyih58nVi5h74HJhydEwDNV6qTii9vkeg
/ktY1j5k3Bbpu3X/lPetuunSfZ6JHlcJNJBR3MrLWsN2FZ6cJ/+pbGXisPb4q1FKyX71DX9ViLIm
ku6k4Ca6v9rlIWWC5TwtzI+xJ2L0eIaoJxK3sp5qTO2sz8QYsMN577zCDXVTEKSPHunswV8umJFO
h6/4v63PTVjGMbkKBDw7ME3cqeJhi61/ZLk5OUu9ajy0I42FILL/FO74rSXXYoGvFpBo2+2lFx+/
CvQRT2XdN6tKiiCcZL+XS1I309tupWhXfAar9UqPO947BBMLWZyZA5xnhoOdWG5juSl+26g5Smy/
hPpbLrfXxbyumK+ZFvYzbDnszBeJl/sH5NWdHGreB2Yyb1etdEqo2TNl5JAUScXlid1LSzc+VPcS
YyLi9TvIqIuIZPHTwM3BnMdtkAJayD6qjxhlKW/DNv8qEfOrLtBNgfAEC6UQYniTzyBrMakneVxr
z6dpqfKz/uhQxDdUxLxmQJbj3+OvqyGNB8VJvfkMqSAdNWt2ig/CCX4od5dp9wj+J6vkHQT1oUuE
8sKXTciO+z3/4GfiaK/YkCliJ8eLJ+Xk74aNZZwnK18ZSPEEK3DR1oPWdhzwlX1jJwSJqLjuCEQ+
ZHcOweFuBzik0MlqPsQTOeFaK2LMfyL4DTm7mFbx0cZhzI4KjM9d2h5EjxwVI7uh/73VtSIVmJz7
Hxd7HYJpp+Aky2gShT2UtXZE8tO7J2snGTHxupYdP0M3CudYzA3/RkufPMckt1W9K263JCCXpTcW
m4+rdme5X7bInbaGkLBKFDX5WKDJgnOwdNz8Rb2UoiuRBVUO7wXwgjaSBL65QPN3hmGYDEItqHCb
LcVcP5oqa8F7AUmSoGJ10dALwubymeelmx9pb9nRhvBdvghbCL3e/byvhqN1fomO+s/Taqd8wJh5
THY/MLsY07lxJZgYYpp+3Gta2s+eIE0DVqiDtCV0xTkIK941RygYae9w9qdJQG+ki+JNdu2LTP/a
TOOq1YoYymeK8O5yn4akBfxsBGAUOR82CsjWd62vlZm6VwGA6/cmaBG5O3zKf3HWD3cI33CbNOU7
twD4JR2oGXs8K2Cc7dvGj+DHIf9kPRW48sj2q40YcqsVovAakk7QM4rAWWlR/Dagfvl3/01B7nOM
OWDJBV4tmXD0FLFhnjlopIO7DMFI18vzkuQJMVhA/yDSAckkzUSo9n7uhAe3187OcZiXa3c6gu6K
kI2dW6zXttN3tT1X8P4vd3CK+7ZU4z2zVNXOeQfLqEtXt/QrzuZlM8NsVElUpy3XGwMi2Ic0R0V9
OG3cXu7HjJy/LkWgqNTeyoxk5zrXPHopPdIieGe1fY3wCz09s6SFfvz98J18F0SQ+77PKPVfGNk0
EUmNyTSqVH0n2WMi2w/laSd9UNWRMx0lmGRqgU1yHFJ13dSvIA9VFF8xRZfW38B4+ti+8DT8fHZJ
guiyChA3COR06O/C3CBEt8Sub8NRSsnxeqpubUJ9pUnmagB5iTIXS4jDX/F/6fh6mm9/x6D8+NNY
I/4sPTUWNSY7QmKerN7DEws7+qIy7J3kzUuolERGGn9ALpSiHjIE4Y+YzY9JV3H8db7XxSA7cEXO
0H/pQW7tl8pGRy+5j5cwZ9r+ol1Uo+weLGZwihEp+ypJ+NbqgcgDu+znzdwOSS0iCks/kMnlzuub
Bt/jDKHHjFwtbSKBWMU4p5e/OIoGhFqHJxX7oGL7hhU1qItk/+YzbzidzkuaheGCSNDg4VC9ILrq
yxt0pbiHZRQqfgpCmzlJrT+8p2huDiktx31jbNfzlj2IH64EI/QSxjEIsq+HMZEf/c534yZHb8nK
/u3DEGn1G57/no7fskWOBTvWNiaJoqsfYIgIvAeMBiQMz47IK3M58jElIPzvk13EDoKaISD/l/2Y
aXnWM04TgT6mB+Qs3OKe63/PdAYGELQxqVFYVzqrQVZxnPl7JW9MbeRf/ad6v31QAllaS1mOE0Gp
8xkPmGbzjrAvldCVOxC+94yLlq18yzGhb0hkdsobAC7wbe3N67jJLhG/oAuhdfCR1LCPgxbify+8
RvosljVzQTM/vgG3mbvRI88WzDYQBs46Mqbx7mwmcUqxfPNv2odHTck+P8ASeC8V+reAJcURqP18
D96FJebau/gS4VQ2dvr/yQ8kMs/g3uMfxay7m4FpTUrPDvPgkNvq89zgulrk4BJi7TBtUopb+t4R
s7yIH3cGJMlc448qS01uOIX1AncB2bubEq7N86UFv6OsnnSKJ30iCVaeOyJrt1uC/iXLo0eLeweu
r/K8dlsPdoFMXAJYQa93YbgFhbwFenh5tlKR0Vnd19oy4V85FhQikOx4OYZBJdjiRIazPPFGRf+I
fcVJoiPk9gr+U/NxX5NAQwV/qIHnxdWHY6Tr/g3jiUZirSk+YoTahqy5F2bvAOZDJUZc8o8Vugpk
zBzG7bE2aEvZKiqoDyRVOUF780Gct0xEuyf8CbcL+pNQVOI+JBbbq4ZTNY6gIO/JnrnbLxqES7uf
E5CEt5Y1SOqgALY0dDWmvM/AqReW/TNmMohHfHMRyBtBUf4/eUQBlaWwI6ns4gdx5A5izuEAFfjH
dAaZ2INpFqtWbL59diaLuoGccUbwnUgAfKImxqKx2oooQ86FwKu0aML+5QbSdSpLmrimEtBL9beF
DTyQUHfHFg27NmLmnRVNwXEhbmtW8uxt0ItjtD7pwjCNxSyZ7YmgK2fDjWlFiCk/C7xbv8jDAfZ8
34gxVFhZy/vwc0snlAIPE+enpOQcKNeJCWNU6Sxf2Qon5R2/97ZbqEZy0vrCyknaUdj1Jh2quSFU
TU2QEvWyO9oJ7iEe1rc2ncSDFWeOhdPbdkH/b4+G1Ra7mkXy/1boPYI92hPQUa9CoVssx76Fo6q0
ZwHgOVScI6YeSTfFbpjujWieL1TZCvC93fln2SoFRlgBxohvc1TzYagTWwN6xhOMUuEaa9yQKI14
CnPjJlOpcPpCizA6TxSzGAPCXPJ6/7ewZnqkpjbARbDvoGHKFfqRwFZ13iIbTfZV5cntE12Oa2oi
AblOlxm0kGJOcd/AZq6J2A5xumfJUhaH/FKrsnPOLcZO0MT7G/NqzYwPcH8KZkZDsoGGA61/an9V
gLm3w1ecUUituTv+zCoEzFIYH14mTl48gjGnnbkdzxj5GH4FPFGGRgHeTLiYxB7MpVEn4BDgLvyg
TSms0axY5aN5CndKtOV2fqSyir9A7qcHxFqNNlpPWJIgFztaTDb63L37og4GYI64DwHzRtwLqT9z
UiGKMBBLj1JzeXuSssudtWkfMGWsX7+HyMJ4PUqkLVFLlUKBk/MtHwBca6bWP69lZ38Twrek6Vqw
vTWENsg9mYjePl013fk7xtMDDIQqyQFGdoXX6Nojat0K8aw3keeShJx5XZx0FH3DhFGL3DZjIBoe
+QSpf4l0CyIPZnfM35xZV8T7j9rPdsGgwV+m/003P7+lgJKJsCGxA+PTtW49NhXKLqSy/hnbE9tt
nxmATYRTaNokqBRaG+ZJ172PboJPT+nzlrc1Af8xw0Ih0NqlcIhIzrOu1W5xr5ePmB4K0zgmVRJW
RvfgeoOk3B4vAHguRwL0Nu7N0L2EngU8J6Zl2p+jDNbVBs8/6LLeX5Y6VIAjfyZiidIzYH40Rne1
/cpexSkC59WXcP8W82LhE7e10v/eQMGVulZ/tYDnWPLiAyK5X/QjZEpNhOdmmuUX6kO5O+TY/sJh
+HgXPHFgMJmJQCIZfkz5qfjztsd50o+v/NWvi8IDQZ/lwRk8bRhyO+xsujkWj/eX0dhNFri3XWpT
ZzqR6BxBpjJt0uUxhCSic8Klb2mOcYjiE3X1GYCSrt0zlC0GI1fLGAuYFSVW9CEZfMK7AG5/VMXh
yR6Ot7CCAliNdg6b4NHFpX676omEa1f+JRKo0p/tEYyzu4wS1g1rKJyk/SfwnkT8uMxneYKy0F6D
pXfB8MsEd2QwrSqFt9xMTsXInXI1oq6fJ6NdzIk9CynUAwqB4dYBMy7UVaGj7cBoKXp08Bm3MDG+
b93sfT106742i6Kcjr6Be5uQJdXI6ClHHzQWWw1W2ZEZeafILJJYRLK1BJ0I5poNgnNgU3gjhDco
f2aMCaWLrV1307efJgJgMKPEoysSlKnPfjkjjznHcPhIrZHuTElA4SjrACGfFqjjGGwsmLp5H3WQ
/Go46MKqr6mB2ZGhqfcvSaMqqJrRkG20K4T/d68qUXGbgPSyv1dTFEZwOotKlhaXfmfuGk+L8Av1
CvyyqSZ9yaswtSEBQFfX1jeoeQ13oRlpoAgi1QKaZwBjfcUkkoE82c43CndxXqNaY9hYpg65QkML
Ww84im6KrMEgkllaOHfWq2lX7CZqIMbFH3VwBDLq4maJxRt/nrfcC/3NCvQykWQHV7vbkRSnqAQC
+S0x9b7WaGLxIfn68LyVPiquhGse0pgbmweG0UF6d2SXQi1WW4fATu/ggLML3pYhrOUcnEh5sYzp
EnSPbnkYK20QQNpeCpBtFp1k5csc7mBTmWuZL9lQleh2l8pvnrplLGwDzuzE5Qbb7ySdpJW+795F
jYtbtqUhCR/no9TDG8YB4FVFR14t3T5jh4ptdsTpK1i0JlgdMru12Wg/7DXQsKYN4ozm1cPN0TNH
JDRD08mb0kwZVhI1EmuNZw8pHCCKJ5kvgaJ0QeFE1vn+yJPEmtiBdopUrQ9cN0nZXxUZPdGX+y24
/tyRuGvMMikcQVxjfLT+LD7urZTyIJCDMIBrqaPoxvGB8kKRnucVm7LzIZN8jUPC+JaRxPiMZjkQ
PdvTzLl2VOqf72nf8vWGRB0YBFSDVFVutAhsRNbqnHK5MOeZR1AdgDGg6iAWG89wJNl119JAQfyS
YvyXcrTXBUseyOOUNnAr9CYMDHTAkaVag8rT2gKlNt1fJNVngFChY2tzcohBZU+RE6+Zcp8l4V8/
KOAdn35C+C9qoB3Y1ATiuGpCbvctbqm5dgduUe0LBOvfW+s6o7emlW9cnwPTCve97xvtVAdfogjR
9RY2NLCXW6F++9BSs+U8saiM1aGT1q1rL6EpyzANli0XR59jJjzOP95dX0aQhp2TrntWSJot2jKl
scD/ZhviJXIe+x8jCKaT0tpFGqZ9Tt0ZhGfP2pFDjTFlbEWvEKX6eBb7RA1MFl7sOFkcEWZvxLvV
7CZipGKIXQsWURHCbmDqudGDRKLwNJU1fUskwRyF85txHj5NbzvzCL2hDDrtket1EGGlwnhUfivG
enP+OiCpGAzE+A3+XgT/PjW4GQYW6iV9JNfD0d6PuH1PNRC0dFQJZqnM70d5C/cFbwy69Iooh+me
7ueP85MJDCXBsG0kJfX2+DTJx7sxqcxfUpCPNAg451BTwFV2ZGTZQA1GQyTMbgdq8fAWLUfW0khA
KJzi7Nqax9z/aQPXTWBnZPE3fE4Bozk3gS1zGc5HOerKLXWNzPcrXbOl1FlY2dZHFEi5w+981OiJ
5hTbOyrpqgwT2DO6DwdVvob7H9VRt7NvzR74o69YSQIksZCVzGVOs1yzg+DpkuH0ckzlVoZ1gUsY
vDxxxuqKCap5XuNZp6b/uyS2mvS+kAWfrAKPnvENG9hzlm8dTWLU6EHLudv4LGsvI6V1oRrr5XTA
9g8gQQ6t/U+zbbsOEPmGcfup/nB2U4nTloJ1ZqbTqPu39k2g6yRCNt4LVG2pSQ2hHXbLK6ir/vru
a64vXTooSEyLOag/CQYreaEEkCiPMKk/UfHkQYE6Aj9BlLscFegzDnMUaunFMyMb9+aj+kiYq/5P
NvZ8XGCSI3bLj1okMw3QaYEQcK4zxSgff9SJSwk+8EQ5MnxrnxpObXOKd3gZmivBxrhD47jHlyCX
n0o8UbK4I6sZCjN2w5V/ranvYheHhs4N1glcoY4/ZJDobIUtHC3ZI/7BcjyW5v48CSsT4cuTHpTH
Wji0cuWw5ki+28FGm03Au/SXp9Omd8e1TFD9+S5oWeUziwWOY9W1NMGLMOi6vaeGr6tJlepBGDnb
v85Y+9FB0gVpmSvQVjKFYKuqeWGBIrpdJhE5ZnanXm4kj3U10e2QFG6kgk5H0cdAqnRAEPyTsO2G
4n5uHrceiJSxFQteR3LRhyyhCBfzmf9bhr1NUeqht9svCEieOFhwr9CBYKdoV4dG7d3Yq74SpuwB
j8rQ+kwpsOfb412HkbFoS/lIJcy6e4wdwRlJM5mCsauWYHEs5ZCHjo3TN6sbO4kLJbw6y/zzoH+J
likQRhib3WGxiwIjYVcM2LoVYjwCjHCJ45FmJ5076P6ksz/hY/PsZ5f1lcipW5vSKBFttNOJxD3r
YXfjHC9LnExxuK427keTPsnoQS730Ukc32MyQ6VAsrSoDuKUtNbJctq4l4X6GUpl5jUE4ZSkhDHa
3MvmHCmehAdufh2/bdgGf5LQGjHkQL68n2BQNyKXHdiLq3NBappjMHiNS76ucJnYl/cboIwqQuau
ILur0gDxWy/o0IGFh5L6aa5a85kWn8Jc/+uX8OEHgBkYy6NK9PZEGaWNM0gTWmqDjNFbK+7889zo
/6eJKXqKXxspyKYdtVKJbf7XcgIW63E5qrzZR1kTVQi5NovchT7TPRSqUfJKnpV/oPCJTDKoznSF
RsOaKy/BPI+/JQHG4epJUiSEpW961Wv6RZMMcMX6SQ3BdJ8VTbhaDzdF2PiWKhfr5YHRB1rzcBV/
4Mf9u0MvzeLgx7HqMLAp3Q3JV4N13R0qJi9dE066XXygvUbaOK8fkjy9eeq8XV580rg86uXTJBrH
Lsg/8JvWrx3CXF1+UEEUhWFpQc+bEMXtXtSwoiNEm740T/pmbNfyyW43MGprmVFq+SxsTE7epVuO
+YXQehD7v5TI8AQYn2oIo6WUSUiHHocDmrtvreM9fMgfdsZBwe2H+3Rp1GtrHsSN90chHvGjOLr2
XddxLPxhzCqbfhTrLz7aFutM3Wx+U/syDIy62dYUS71+N6OseulH/lXIhh4+baDOfwK7Mbde0mSO
O3Ld/gd/beDRubSoeODcW68ZgpB+R+fOoxLtCbevdgGgGh8hkJCnaD6l6+5VOjV99XsoZjQvhhYk
yG4F3Ia5P34c9lHSTcF3GASWsNK72uFdZaWNsNTyCKOmPrcOcM3ZaOL+bR3o+naEQ9Bu6aKAtZWg
8nJlSKh6Hyc/vwPcNks2PBnWBwP9havM0WEZy/5SoFdjb8GvUx68pLoPZ0PTrw2LJuKCHJ9UtLno
VqqIfBqSIn24EohNLmHV+LEmU78/Bwgkmgg/LPll4KCHDGk0BRXZxvwe2HTB36wN5Mo/pEUiboTh
B47rtH4Zqviiy8D+M1mMxHjZ9Q7OHedTsrfQPwCGpAa1FUOkMBTtWBbKp6Ix3S9JjMsAKj50lo0B
Gs5HhZjOjmvfI6/TW7qJZieJ1rSIzafmJo8pSIAtoDs7GnHKENET4KImxUXEIUUasBUbaIxX+0o2
FcJ/nbVsg/XRbSnAk0kluUsqkEu/q0qsgK0zsSW267BXPeL0Hq7NFru27KkY9B4jAsoGzk1AT1JO
dCqtWHz8nRoQnVOV5EwnxBS3dHvUqy0xcFCi0kKi2VRLA72FjX9Jko9KbdYkmCABHl+mzon+l2Xa
wD2Gcc6RJ4dk+tJbLxQSah0v97+lTLRBmVtll2V1xAyj1kwHi3VJifZ1ZG6J0k8TbKtlDNbMvqjp
ux+kfCxAEZoV1fE/48khyB/IieFMIZN5nNV/ze3e6PLo1GSRNBDcWX4HeVJgknVAPW9Ac3cq3mhJ
sEwvG19ohQMEcxo19L8f9nbIsz85r3ifeS3gmcqI8FNsQXUN03ftRgkiuu5gAhSCL1CH75MGd/vk
Uts/FBHVHKW01psGE4mSg2jYuPaG2Wg3ZXq115E6FcSGha6mcQcLtksPBbx1S26aV8/ZwJS/jIBG
OHprWnQn/dIqd3VSlkRgu2qNGFr/BOQzlDnP607U+EOfZskoAziraLtydVEGEpHLmXfCDhoQxccB
valKoJMYQ2WipKgnkaDN5PEmHcMdfvazN/MZX0XHT7/ku2BHsTwiH7ePN/xjPprbIqkQGZFjkSjq
z2utORVQobwk9fAjkITC7Y93Gp+4Hlqx0Q+x9CZYTnZ/+I6PSwzB/Xr00NvzIHpeZjtSbqwqwgZ4
pTX0ktkLTYq8Zc9bt4HjnS10JQxwQU9dV+Z3HgsVU5sTK2c/szn/FKS85SfEn2LwUZ8h4iJxs5FM
02tvNthmus80PjYF+4cUVwj8eOQCwpMt0j5nKUxcC3OdHkYQcQfAk1KLKoBKvs7eQgq2rg1Vsgii
NVdOr66yvIqj7A+j06NO+cwY7LIehEh5kfE3dAEjylp1sSsfREmj7BckupCnjBzK05vLbuPdd046
OOEW947aoQ070djpeJjfvGCSdA82YwJW9lNByvxfVGvzGBhB9lUyhjOEPYrysbpv1pdAneyWCg4O
iPBuUlVoaDcC0gPtekG3pV8HixM8n9nZKkglcOg+s2B3OBwiZTTc2EesXNlTqrx4dHy94giXzG+j
mcBaOaIu6UF7priEDOjTjUeDHLflnsnJkiA8AXMK3Kc2HfzQLpAnuZtQffW/usT6Gpb/GtHVI/1c
E92SchX8u9NtO568eMfEO9R/UmGxXlrJnLaOP3ftcES7ukMQwE9tIO3JsIwQfFtGq+uLlAPINHZY
qxsEUdoPIoZ/KvSW9uYPBBEBTgVKpg8i3UCgBNqSExdXJpI7LiXDsa9JIsFlc6XVskq07nvUtBUS
tROpWZgxc0vynjFNyeimoDZB3TixUBdDLEXXoiIir41BHnAi+vlToi3yEc4rhWu/ikzabcYzinJ7
Q4CQbZJ/dHnaB1yku0gd+girtwBJUZfqdGNwKJYKy45qcw96LIt1jh1/n8peCaUikcKfyJ4lIhy0
dGKVYF7KZ7ackBbWsf2tuPDyCmYRJTVCPZS/DhYcWbzD4YhgH/56hoGQ1Q32QRnnYED+/4clNwdc
DHeSwPfC0VWVbszQzqzvjmnkrdyHeZn3XGIbcCuXwiuMaDaktpM2LtD49TYUalaYUG/LwQdFeUF9
je5Y8mh1Zj8cQPc870bIMUUWFnfjnrAzaKc+NiVL5nsUkQOUBivkYA2RQy3i2n+KEvZzLJikkZMk
ytZp07d6L2eoQ8DxS4ACyl6Q0Za1pBzx24TNkagxMFBALXCR3ovPQc4FEmBAz/mVyCYcTLUlV59L
7kpvbBaK9v0Obla9rt/jL1iqbcw5PaeDnc7DlXQJpGWWGNv9QR29glFICVfvTBfCiwncE8mB0WkJ
bqAZIqJ70+SbM9mEVlOB80foS40AXH8C35e45dvvZi3H8nfxMmd1hJZ/vkVb44ilvfQ4Lnnuu1j1
27RseXUY1UcoS7VR4QZpwkHUqePDRxiz26vq6eyuu36jI1zXZskFy/m/Eb9jLha7eewq1VobGNFZ
ICG76cOOjJR0vce+KU6Tv/UbovJYVMVKyuwJCnw3kgjVXjEMmbCBcNnuDK19XuE2xguWmRuetOLT
1WfuoYOo2PyIAmW5gthcNSszaCkUrzoVk33KDKepcTFdqfsPaDXvnRhSxHn2mp2AOYfxGcitNM53
2C+duBySP9Hs4zplz4vozzAfUCs7monAxkGEBQKqaLd8oyggJvtl1RMTDnq+0GwWw+qF4R8qSOcI
RlCQErLAb0uNQhu0RuOIsysT9JoWtby/oWOlr+m83mvOi6PR4ATeiISIAd0X6QjG23ZddFjiVRoZ
YVo1dO1KJhIm/hsquu2f6t9P5me8tDg639qs+STbPsAGhtLBAc8vhBwPVX4tcDGs1RMQuFpm2128
2rPeH3Trfp0ZhViywdVlXvhKnPI5+Icsdpj1XEsczRpIzPP194oye5C73RqDxuYSD4+RzSbEuGFy
cDgyryXDvf2EdlPbjYXfLUjrTc+3aZ0EJHiVGNCuESaPI+OtfTMykdd+3xXD/hTIbQkjmp4qoN71
gFILbuVNEs7qV7TGCm2LtzWwlO45y2yhW1Qtcc1+tbyHrvKlwWd8Irb1o4smg5G8JnC172t1CjOI
2JM1aoZOiZMUo1eQOM1TmPQB2J4kXlVhfLpnuZB5vCYDKOr34eSUqE/RENKpw/Ehlj5UbhY/231a
rOgq7EQHRQOwaHxCv+n/xOY3bPETMMipaYQVrjic1KvqMy2pmsgVAKl5OePtFGAuapG3I2/scT5f
+KtHxrMuViITAGfnZ2FHusqlxsyKgmZoHjcWaxElJ1m7cxyZeDbPCMQVgKS9spkkAh1y1uFxrH0M
4CP5GOhcKTWXv+vIzKzBP68/tUfFdYNSfTM3z72aloMxHCqIqLZhSYl4yHI78Jwr//2hBK1CAcHo
dFqopRvT6m2dXL1w6cBojyNShj6+2JMK6+luYO+YGN9Z9y+EeOP3Zn8pgEc+CC6drtdr4Ep7ZB53
DmuVezatQYbsIGSR2Cxkgb04BNbWWBh+L+uKX7a/x3MlFTJ9s1tX1hAfACV4E4zHp9ZXPJWKORVC
HSGd5/541amYwKG9e6L0UCFDHZu999k7oB1GVW7eqsljkZpqzIz3uCWqdz0JtPvjpMwuLzPb4rJT
62sknDwqiMFpUEsTkTEwEPNFh7EcjWH1uplQbem9OeuIQWfC+Fup7tZMguGj4ReHLawv0Qrduc/e
+pfrcf/xrl59Hxa1AOH7pOqp8h4qSSExFKNIGIJMKgQaLZesn1nYrvROL3i3aNDKXjwLv1v4MYXp
kKzdIlU0FdFTC8Z9oDb7/jDaDGor9cy4F6iorgiy/EhU0VP+F5eAsLfZFxwKiisrow09iuhwxrlM
4Y+XNDuYAM7Hn0Bx+lYVtp+KnYyf1zZIGdFtyFyTktwVJbAPbIikb2SlMr32UcH8ybRvHvC8QIWM
iH5MbK4ExLjijpaAAPFWH7BZGdvYFoH9JWyTB+K7gbX3XMB4Ghw8D664aPejiwZpyu1aQxj9nrXP
Aay5zcKwL77UPL9XXE0O6S5EutVHyLGtc563xgvF+XhIpVOwY+wtAR1XomgTjc65x5aSFfd3YlAf
a1xhIvFlMNVVFMoet3e3WIGfVmgCEPKp5arWS/B/a7Yj7p/Uaeot7pSl5GhbMgJ9sTli+bWouhdz
IELyxp0MuczYHtd5CrjWZdpc27imSJn21kslppQ/dMgVYUYCqzCQyAvpTTXQNiDSdwgxpmwI3zF1
flgSUupCf46ftX/Lct8ekFSw4uI3zeC3i+lOLJoPyMm+iocGDdFJGNwNIMl/xGp71ol072hcZe3k
K6yYGtHQtXyxh3SmDUBkouGLRTMz7trr5fw1qUz4DxRzwykY2tfVIEzNHR8VRp6R0FNX3XgZg649
o27lZ7lCiCQgG+Q70B3ddw65P2kUni5a3akUggBO7DklC+m4Sebpz5etUCk88f0VfmdUSPTwPQxM
fD1SLE/EsyTJ4q+QlyTfciozmQ9KSBBl1IpVSSVywQxPWpp7jGmz2Kp7Kfl44jT3KFJqjooU8+BB
tQgYzz7O1fswJUvQ8h4AKzUdV/gFl9pyTh864ASEkSlf0NbRMLbDVAROtrXC0EAX2G6QhBRMssCh
a3MMxnoguzdL3vSLN3ZyzaV2QuasHcX7/YTNZgG2nYYBhNEhAGIH9gxn3htqnw1U4hm2g1psnH8F
VTF3s9bgCT+2+SKJNKvNXCjAlEnRkH68T07z30R2+yqwkA5s6rDLIkp0qnpI0VxSvm2HfrDf1iIG
d4p1BlA9iz15Qh6IntadUqrp8EklMIaKnZrldPaoRvie1CeBs05801HAE5aaFC3rPdOR1kjX4gwY
RaY+BgdVbG3DRr11ePj2uOqWZ9MmsEiH82stmOaDzXXbGHt3b0Qk/UjmE009pGLEkRHpJ0k4qctB
733n6L3YZ1ILw+VcILqZjj817XAw5/IN88IqCOReagsCCMt99tIvlQBrKm5ThhaZkFggop+aNQz0
0p/Rr5NdBnIA8T0Yg8dQ1J78h4FRECFDubbLN/pi9JrYCn8zv50JE02K7MbTrl0bjMRw94+FkOKk
5C7QG7kde6XynoOZ+k0NBpK8VdH0osZn5vOm69wxbubvKTXpwG/w2eCS5U8aa1ZFgpm79lqbW0NQ
y3/3udDgoHpRsIE+gI63UjKxi+OsK4PO3J1bKDQmK3m7NMjp8vtSVkE2fcR7yeRS4NKKaToLjJyd
wglGYN6khHZFmXKrTDyW4QIMlS70Y3xk1l5gJhWvsSlSWpN0AbSdj3Xs5QLaT9fHdNTvWG/sfIg9
xJQ8R8u6h21Esnwr7t0IT/XHlxQa23PdUm5/2tuxK5QU3eNp74cj3pDTZnLRYYIUy3ZaUz9J4JhP
nUHXpyacYI1S8fgOeKUHBVoLu9ZYpYfJ4CH8Y1S/p3l3cWOeON3ygVeivbBem6Uv0ZnlCRuWJy9m
2Sz/DIX31mPuh5eSzHSTa/kNpG+a6Qh6s1tQ9tUTG9I2hmqEQSLg/7qn6lUiwGkqbwZWbHPID7Yk
XZwREnxZM1TVQvaPfhawgMBjaQ7Tvh5cT2/OPQC/xRRESAPHIs3qUEaf1JVEABXjLCDHf2ew43vm
SDZZ1w2ntTsCEEFF15Lzg3NbdgWQzQepVg9PhlAnw8IeVzHdhb+tFrC+NBBJQBNZltwgseWX21Nz
wSfodZfUsIzufH7yE9X+4rEixOe+q4hCAMDZC0ki2YHQ1OasreneeTaCWa85sgHTN8Rn8Qjm1mvM
dRpXfNg3TSU4lW+QlIaQOK2g1PEmtUXrP3hTFTgXYh2INb0HisyaVIN74NCd4MpfF9I5zJZe17Op
VHVofnvdebjwGUmzaiuxiscXr1zCE7v4x5MqubJvx9XgfdLlPncb8+5Dck0bj/s37rq2bqZa4gmR
6tfsL+bm1XyJslcVufXr8Cib/2nL6W+3LLoTdIxWmKhEibWjYFDb4HJuPypRVPIYxBFnwSg/m62j
vUMwdWlx8r5ociWMf7yF/Ijxg4ZzsF5t7RD84aFklUupYM0DV+WRA3nTWM0JKbT0aj+/mt2JwYWX
2zSDPxhK+7PNhH/C8lAaf2lbUnz9u1CZBhJtzgDK2f7mw2WSArRaks7S6+j+v7ACn4I9VXNZb2Wr
Ntb7I/AL9wrXGPsaaQjye9pntTkO1cb6wvYMSa4Xa57EcRy3SJ2hxGqzhNx+ED4124WPjklcvl+B
uqlwXjF6Znixlg7uKpiXKSjflBaYvq6idekGwMbvGtdxoIiXJuLcWXJqESAPybf5Pzu9ZymCSKAW
KAjxHH/X1chvQUaEysVek6pnWwuiNCM7GvwXgVYZCmrrI5J8zJnmPPGlhqTBJmgCHAHicW/TNY6N
iJsxm2XTt5vXdG4+gcvEtGOZDa+zpw2B6c+qA7FFSajDQDnx9mVv+A6vJeqxuhLK71sGZPUhNZWT
V7wMT7yvRFEpvCYW1EgTuCEg3UIXqF5+jwFk00+quIDc0PsTuNijZmUg1vJg9wi7Dsx+ywdLbjEA
jiyybLM//zxUNWkRLlIm53yRsMblrSdjhffxEsqMPn3jx3w2c6HNb6TDZJMys4GFRVUnxdir6UNV
JqV2cVDNplc6M9lxc24UVfDIbrg0r6C1GOe+Vjrt4GQ0N9tyVJM0KDeohteMf09dN0Zq+OznWHYD
Ij2eb7iIQgxU6cWRqM/otaKufiiJsqab0SpL9lPoHVmfvWJeRq+yCQ61x454k/q3tjBr/e+nZ+s5
iZXwmqGDgKOOLHR2zObA+GwoxCvcjZiAnMq2V9Z9H3BlNrmQrMbS3i9luPkDpsk00CgifohfaceF
eu+tXW4KGhsr/IWfcOeAKkvJAY6BnxhtjID35spXJw8je/xqqA3+Z8p3q2UYICibpnnogm5AIY7Y
vJ7ed3lBhfFJ29PDww3t1Zsj/9omZ1dlrYYq6DpJ3ePCO7uayrABVYGoUDHSKoIQPdfp26qOepO6
WM6raoPRtB6E3dvTlNVeaci7dhHBFbQh1whPrIlLdOe4ucxroWQTfptGt31fl2drtdt2Gkj7zml7
qQ6XE9ubzAXNTmYACzySuLcfxmaDhuf9U+n9rzOfju8DHkrEHw8rF2JCwDf7U3Elrbm1OazYZwZv
OnOFNjFQ/8vzhR9g/4bctg0FxFNEpHBliRitB/lkNoC0CYlUzMBOVxpklaoIq8yracMwQhBNQsty
QcST+iXYd76v7+4UWcToKm8rxwUeWJrdShmbwQ5CeiwRoETAsMTEfrhWZG536NTJL2yldUzU2Q5f
pOnE4hEE6wrN+tcouBccwj5cazT805VjVMFpqxg79CQU8HnOn7S0Z0QdR255CN+5s/1y9MzlCmAi
pb1IW4Ak/u+tX3F6S5IhKgAyT13+4upgqaISPu31tBZQki+RO/DZS+FpeRHPiWsluXfI/s8xBzz/
/O7CRGx1oudscwlcwKMAW0X1JB7zUnlKRyfOPKjqj94diDoRgoLnvruYS37efa+012Jq2tupU9XT
ZKaZhQPLfTeyTBD8W6cXggkv0B7OA2q2YKsKOFv0o/X9/nPFqzKg4IOW1tR1xYjizzrBh4+R3swt
oaz5ejoi4o48lAcueP40QSlRyQMS+jW+lmxuvcK/2Vc7L7gP1cu6BFwI8sevsb/W64MQrRNFiOnx
rmc/dKKfqTY+CYz3FgF+C3x93ttMrsBzLRMXw0WSTvB7vFrZEFVl+mTfhEnSIE3QOkgTxi6AVsF3
ykVH6z99YuMtaQUI1Cwth5Levv+UWLTGZ7Ol+bRrlZBTak2RwQipiGembzm+TddKmzK7JlEXPtXm
/tyfZbVM6FU9A7VQvqQhxXPr7DYNAKCeBEB/dvnuJm8C1LUvfDeBko4OvC28a06sk+377BguelaE
tC60CkF8SH6CdKwdUVyT/aOidHgYdCdsjmsmLNHBsYLP6k2TId93mVzHW71YFiIRgl37z/zSvspK
0gmMxHcifxmXfpgYvIb6g0zXAbcnhSHaCa7s72C7BVIFzCIRWqLnr7ipzHTWYHNfl57hx4kFwDJC
2AlH/MmNeevjeQ285IOoMZ34h2tGcWx/QTELC0dG1mb6LQllijPPpIfr/wxIxI4Pw04INhN7L4a9
4fFEicVrFmbKmiLDHB88xIfZ4AROamz9KZnUztPjc/oLQHJ9H9koth6FkrUyAPmigf2OIcfNkiVt
k8RnAcUcFem8W4kkadVOvr99gWJOoD8QewYgwvQLBypXZ1GZ3E5X0p45m1W8iM/jlw7W0ggT5hCs
7tTNsynFBaHSiDcmRWPyF4aRSFZ8ju+q5SAWlaKN8OpgtMMKjiMBFZwMCSo5giyQM+4oLsICSGdY
3Cz37xhlZJeq+jbcgkArNNFBMooakm4G+NgJVs+alfVS76+faKCo1DKzpkXa/21F/CgGp0RV500I
wWaDh3onBfI/wsFc+GuNf8AAayUYaOR/600Xi89ON3bPL8BWks5yZpna8mkADIdJVzPm32uPTjhj
WuB7fKgjO9cRnniHL3yaiSHzKZHlAcw4XlXr9dJDngqL9PRS/OYwlTPXK4vlEC7wOhpLnUQ6kwy2
Vs3Usshpn/0iX4mjK+ZgJWITyOifoiN/KFUuHVXILJhuT8uM33KZFOMRZJcz75/QckObdUwXhTgt
ZtqKbQJHe7oPcyIyk4na62HRFjQ6NdxEMu0avgeKPoTpWj1gCWUeKtu+uh24l6qnM0+txTPmf8zu
TDcbXiIfVd66bQkJ4i8yCwCGuAS4sAuCFedhbmClxhstVlwEAcpwI3wqbyOuMXX7iOB6baZNv+Qk
5TA9uLuN2+MnS2KtQJCS/9xT/ip1OHpxrtiYew2vbjapDoCvgqRrvtSjhaZxQSH0DPz1+cuP9sEe
eUoLJCdbJhsURUIgTmTYww9zhONSLQRvrV3zbI567s0kkZyn996IpVtouo9WYtJfnc24sNNSbV42
Nz6p1kJF1I0yPb8/p7hIxIA4J7O0BryOiO1/W9hRib4lb9xNB4YuYUE4ux5OSTqO37m4ebU22Cfj
h2zj8V4opTRdh/54rw8XFBliG4E5yTC6XkvTkilMFX60bwBZmD2wMsAYBGKMxE+Klj4ZtVQjSajP
GE5OfbHg0SzJAzHmG2ZAinsXUX/HZk5wyMwly8x+YINs24A4Z0N+RigCW8gjuTOC9Bg0KsUmqzgk
DYUYfzyAV98cQA2XKVupxRgXLK5KKEuEPiDE9lmM2gATFNVKsuldmMdRmw5gALGxCg5OjOAS0x1i
ejnTE//2WI6UmKMnynKMU/QJaZTovf/WOcq8AkJJ00upsBfjKmzDjyimN2cTS2Eo60rXy9fH0UMO
ZbwKqIvNSKNCLVoGOaFvP/ZcdvR0JbWuPecgs1Qj3C05Tjvgs553RRwe3aQUXLV81aaLc/9ackhY
o9zKPksb4yYdzHlD2Yl6i/Jt9o6uMbaJpDycng4y05VRcKeq+om0YMFhttXgOuw3Ip0F/zP62pQS
rw/wxRRmX5WrI/nZM6yul0603Kg5HvZs3KWe2mSZOaBppfxX2RZqYJv2ykg6kWcI5FRbbn6lI5EB
Gb05/7S23Io6OLKEaJgULnE0r1Rf2FayS7PlwdIOCyLG6meJzDJaAN/K8pObpZBq3EEp1oKrqpYB
TTLXxgjFh4JW4wGpVpwdMxyYWwHgp6uoruRIxVbE8lqAOuDXgh5Nu9IRsQ4P7DzvVTBmXmMtLxQq
/RpYgBVmTJmpsvcfT6NY+j3GmUSJhkuePD/lYoiK8b65mgVh2z2QZgg9N9NgM2Yr7NtAr5bsxTRt
0r18R6sySb1mmfrVL9pklMgY0pWNivnLENZXtMG8mhnyER7hyQUglHYS5BB79Qf/e7wMYJOnK5ND
OmiQxN0fHY1DXzYYM8pMEcnRBbnnO0jMiBoOoXeC+zbbwEfelHpXWfDdGTG0qzyxpZgWxLPfgf7j
oJDFgc8CWfPJpeJ9rP0y2XGrpsc1VVGqV6t/fnzlAZfUsnzyTejeBkiQcpoXMGj+IZXRsPA49K/0
je3MmxwoeDtXhbTEdlogeCtwmozWiQd9T0y8wzrEE6EIwQLJMmQCG2NNpXTmxHRSMKeEJRs3wu4g
/y2HZYuNtgsn/w32pGnTecvxKC0DrZko7e7LfqaKZoFDE/FFRpU25x3xF3EqarIE5yZU3FFoiNXw
/DRjIJonUzYgsmggFWkXdbycHluyKAXoLbdlM2WWB3LXZxpaHovJtDv2o258sV3Gj15UBlR4PcI3
dbu5QSHmXGCkeXxewpHmtCNI0zDdEgkpjlKh/jiku6gGQncK3L1JmVqLoGZwje4UWFQpzS0y7e9O
n4sVfW7FsRKklKghydIOn7RqULyUcD6fwyeKVQeAuUR7pL410bfzv9DAGNfHdUQON6KmlmUUBHfG
wkN5YSFAB46EpjABz5Ibyot7VTZmvGfkqSEWXvSKljjC30y4tRXOgWfQy76Ejt9maAfFkIlVabAh
HLAgD0nWzny/NEd/Jp5KMPLp1UPOTsAf1SJf491ntDfm3tIVpnX8AoFSFFnqx0v+WQjUUUH7GHJK
nZfcZw5BZSub/4Fis6U1eTCtaaREvnoqUvmeXgL004psqfnoC8lBrrVAzJAdDckgU4htV8WnV/Hd
kBjajLY3N8ubjCT4XfJacSyj6p5J04665gyGbSiiJdJNGhG5zeyyRQkw/F647G0tLbMPf+NSR+rm
aoHpHxp4BJcZTvt9LqPjn+etHlZB9cXxwEzgDL1VI9W+U/vpkNsRLP66+uP4Xic6nNt/LiR+iYle
q3D4YBswyvOuJcneAII+zO10YXQI8koUccncJqf7IDHqu4F6rtrKz8SRI2Dk+VXJL6RiH0oq2vmS
6+XSqUP/JbA32VKNXQjcbcUzdanu6wNGwdZRhsRP92LuxGomaoZZAMVO2VBDtBX30sRyCpW6OhfH
fvFeHfmZ7MByOWEGToOP5SRMhbd1GR/IasuXtVzSG1EZfJ3i2f3ZQSdaMuV+ChZ6tSLfYd7n6c0L
uGy23Zv39y27Ax8u2Ktg2tna/U/Le8t8o5cJx0GPBOHAm13QqOC6lsLiyITX2hP/r1uDIonZd/T1
37WCVO7vC0j9FF0KYI7yTy10oCrn4OR2Eg2fWP5P+uDW7tJQaHFxNg3gwJCWOCq8hJCc+nEyjEsK
v5zGhJ0HM4kNBENL8eLc4yj5MYDh9RgwCyAF1DGj+KXnCgLqeXjKJWuo08FjUn83yOYsnNHu55Vb
ugKal/TNWEjLCpHDzggs+N6DkTIa+1/o3Mg1u3BdcDYCDAM6DcsPjOQyYUzvK/wcmyqtuoze3I0h
MeiC17nJpXG+2bBpkyY3dzGg2vHoZeN9AXsyiYSzajCc/LZbA4E8yejSQ7IfuQgehj8r7VMTWvV1
rZNOfKkYhc5rw9Phc2UwKea5lh4tym0r1N3d2g31XNI4Xzw4sqTlBE/pXKyctATo0lTDOpEWVIYX
5MxDZo2dCBQZ4RnvM9xozEhRKVT/Rbd6/2Vk7UTkO25S8cfqrZzWagzLSFALbEwJ3qIcbfj56KoJ
j/5nO24ay12LJot10z2bBafVx3ZHSqQ8PtVXBeETIstaHty4scKr7oy1qEJ+IKufAuGx94exaSau
Elr7ChG6Gl4ZxZziHBzMCPUzo4r0SspKbYdFFE25Klrq3UE9GRMK5ve58pFHtJsGKbSbLq/MgsF6
I6mLzBIsbqPil7vPVHEurRxEz18fK1ZUoB43uEK3uvPwoXwUuZZSQfbn7nZZGFy+SeuqmMY6xHDa
H8LgmoRS0a8Gkr3p0s3eMIKUFYhIp18iDRxt1ajgBnvRNTlnh2t9e33rGYuyBBA9X8y2wpOpGU1G
TgWdQQtMsSvWJY+zMYiGcxVfgWmB2BF6gyb/2iprfLUKobtsAgrVkHBC1bFPckupalGSxDYw9JCP
pr0NfkTZsuy7m7fCQdJyUdRieWqW42asvJy9ErzSEzbu/oKZjUSoOuflq4DEiGee+9ceVg087eVh
x4Rv6LN6W15kqnmH/cFg1fejs00/INvUVTs4fvM8WJx92I5W6VltcrVGt8+Y34Y3zJp9tTc+qsMJ
oBTgjRo+iODEd8IVYWjPdBge79+K9dIMSumy5aIlJiZNFxSXjGfJvYIFptkry0Dtgt5+oetzE3Ry
Yck5X1EwS/YJjwitwaRx+pnIKZXEF3uwfE3SpYRdZThwOuJrQZew4VV7Grzfuqa5EEKROwNc6thx
tt5ply459A4rD+Y5702pW0eVMR42h74EWm3huh15UD+b1BB+b6je+8honNzu/jPpgpvwSEoH5S39
cfHQ5cvK9YYEDn1kXu5dgO0NnxkLeT5hrOy8dFQBQCH0NfkAqSEmXlcWAl6CByd7zRgbIIyZiDkG
59e4EXVJojCVfKI2jrmmlsXrrBl4vWhzGSgHhzmQdVoV1B06UQftqNjBrdDUWQhLFa0oBkKdZh4z
bKxzt3CcQajRYqxREXwZbOO1izKqJx3voVvcOBhnDyWkfKK92LWLFxH6ceZwwyjWFRIQ5bGkMKHB
+bJLsBWcKW+dAYI4c8tyv2tPpiJAq4NRzuO2RgmqEA6kl5jHoMG5cX9UDnvXZc6TruPDE0OJmYpf
WAJcyNtmYTVwnGPQtu5c7ZUZDQkJyQ3Xc91VdjBUOvvCXEoUY09RifIWqUHoI7olC5F8K2wAKZlS
2sxJPmP2SN6dH4l7l2Ai3D1thsV8V6m8H2so3PJ2JgQDm+0MIGKVOgOV+jr9szvmuZhLiglIXQ6Z
Hb+BwilE/GE56zHP4lEM5R4oAuZYZL/lhuUJjnZKe8IGDnxiLAJJEN7saqW0WM4VK+CvgbE9q5Ol
jZlv3SPwzAZjlmNSTdSNhelxGHP5E8C8C3gNC93SQ+qCsX6KnM7ZazwHmJlvmqPbLYmL52n2GMYu
UcJT/rNJfZrXDp73g1IojdWENrTK2aQz60dgK1nnstTPA0BdO28MN7wcuX2Rt9uxeAZUA7/n+ZLq
zyDPH9a1wswBaN/rQUXeMZ94qLOQ5R6oMTqcUHaSsO7PADDm35ycOXOBPU6B0QzlZodJfugyib0P
uH6cwA2xzU5oqBZqG8Jrl09F4SHoFA81lXmHbIg5DGJsVgtjeNlCvV8kPJs8gfDR0fxe6N7evxZV
VGuBWu3hy57mJUpS49h7Pj4IsZxVZykYzzCB1M9hbM3HpMj2Jw2w9NpTlSkbOdD3FfZHbeaMsGiy
nzN0sCPxAClsTjPX9yAILStnxGkMZ3ApMpCJyGMHTymg6lEMMCilyh4rxMRcRvHM0BLM7F6vstzN
SJLM7SpE2izNhS5f56Od2SzNMm2Lr2MhTh9WfTcI69+SGLtT0spvvd3UtMI23HxRKIg3y0vSFhh/
qy6Y2qshvPxK7jv4jebc2YIPuzQVqq89KboWzlf42rf5RuRtvS2nNLtnmpZGXE8svgchrs2e8YZO
uFGxzJUGgcXz8gJl+Qh2lyLvqWyq4KGnZMAkkWkHSX7YordTJimWhFcB8HG3TaTx/x0QFscJGGQm
9UNIHHmEF84liaQHG+V8ouDC5JoKbWxIPgxXyieQjFdl7hz5J+tQapiDfycEpIeV4gzRA4GHc9Hm
EfJYOgoCTLjKiMCA4FUsyAJ/mgq28h6OwSEOHlgTY/JpSzL7z6d6GR9ouX8Qv3Kxo9EARlrV1vER
yFNz95OJyEFT3CXd2/yBpGjt2KHYVy5rD009/XxqxdDuFJHgB3rg+kPCH4AaLo39q9j6nXe3Bxun
0Ob5Kd2vWFqySvsXXj+Wd55xt+fsdW/L12QLRFtenJ8fYjKhEJI4CVUsKUzRrZ49uh9ZQAPsPXaQ
rkIdO0t9ULIOvSF11qa7HzW1OeEnXXz10p8ct1kd3yiSW1dCa6F06uMrVEHzOnQ8w4UGPDDgPoOM
VJXzuLaEsCPHWTDjNgmh4Lke3ZkzwAVjpr2jTXm/YaslmFiFsvJ+KCaTB0/F8tl+qOWguZS5kwff
PKnJI2TTv0Lvp1JcGr1AtJHvDIGKHvZgQVwEobCVLoW9oW/4q2dVLN9DnsGJWSnBoFBGim+dIWQG
YPoVepubWvJRoQbWrBu4dIrLSDCsveUK18pU1mxs+Wpa6nnqWswYrT6JjR5gVDk5cpAl7zv6+Eov
dnNuOv5+ntQiiVfahSNh+sqc1AvI2se84ruPJJ+9uJjO/pkXDjksr2MLFo3xB1Yuysb3cDBDut6W
3tAEtYi/2o2ExBa3NnhSvgf/wPD5rnk7H8Q68ioEpljYi4Fv+AFyZIa8MWjGKmktm7IWEnIhx7Lk
kEiq14zu3LCqk8zU3i/N+ibI3ERZ02wsIJ3tsMiVFdvo2yqPucOSN+y09ZWUL5jyxnJ7sRjWdS0f
gVhshVYbldphcthJMgXbl1U+Sn+CTnFufBbWOOpfHPAxiPS9XO4isKZKYHvtbKig87iWz29kVZVY
7XKLaoRLIdveoc/kC9m3Z6PGM1aF+YLHMSMTCiSNuSQ0NerMYQN5F/2W3CwcxwQiPhP2F2cJFjvM
Z6zU9vNBY7CpJzHEgDfBASFipfzxskVDw4T61EmKV2+SWXmdqYsgJWSBcJO32641SK2R/IszGzrP
j14HHuN+sM3+BiU14VyMYeOvyhUKokguBI+TtsOYuL5VaX87Vl2jyIzwXOGO1zoZv1A3Wg3ysRvX
QS3sxk+xbUQNrK7qfDxWU08ajPN3KQrlxi/+MBW4ZpTfW1o0q4lkZZQfETtGJGdc3TakWMhFgpj7
MrINrdgPIWx/Y/Mk92zmYyVHJo2oYKn1oetVRhpwZ1wP1e7EiQwVKi4zP8j86NAFQp3aixma2TIA
h3L670xvKZbbWkut5ymEkzqDXNXiks4DAnpmIBjC82STLLx8EBCLdJfnloYW/h4y6Q5i749moSlo
xg9GObX86EvP0+oY1BrpTK5aesi+wjxHJkYzVvrUc2B4LVlu/ZypWXs9lHGrLEDM/cSWD7mEMw+L
8ShF720TcUo5d9XcqomM1GJ+dY6pr9IEK8E9y0pxO20GefK9ehxPsDrlAy/8DALbWMYvLyPc9Syn
KAu1xubZ0UsEzFA9cLPQulkzfCSHuoVWZt0Oy9n86fWUezhsncMnb560HxHSTHIq4wlejNRpC+Tl
zE7APUvf1JqfJHysTf9H/TpXa7aN90qjbVDz1IzX2s0SnDGrM7HrUdLVCDv6D+vlmfcM94gs7ezt
DihRmctyeNXtXtvfTdCuW0JgDJr0s7MpF5ZQ7/nId2sFMO+S6ftE7FzbW62lbun3nnJiYKDXb9wF
SH/Htmc2LztTbN81N2N9/FcFwzvPiCEwhpJIpKMUHoaknXTVCNZp6/W0zMFOo3nglOfLjbyGx2vi
f8oAYNIXPP4s43uujeBv22mcHM7CPM3Wpop2vLOPgqhLlp40GyslnEOkVjbMgVdX57AT842WPyn/
U1Y+il9LmcbGO5VPk15PniaBjGKUFhX2Z19371DXlSlgabASiPyoIsENsGT3o6OyRTDKd4T4xGfB
TLm7W0z0bAP/cTAUNRX3znPTmM9Vrx5IuqHz/89DmlcssZ0zab+qKMuLlp13+iXrHzb00Zt8MGGl
WpQab5sVTnRvTyQo/rgig6QkQEDP3yBx+jbXeoMZox1wdtAD1IYLrXBNMEsIQuY7IH33Ov1SqJra
+JisXDCe3ljHXOeEfy6cjT9gxfTmsse/Ecfj3KWZ5MlOE1Rn2vlPKw2pskiUd0RzQ8IgWHGZhKLY
YbAyknpU8T49qZ+TJ3fjdvKF4ZOfUtbyQdhqFOhJngtekCOz3PUm0GYjuKTqEiDqJisyk52+ZZaB
s5wwwKa0wmhRIpy0SoEoAqen5gIsz9uWhlwDvmNdcF6QFsiIUT6JNqxPUnRe7FlHC/Rkd7OqQAwt
YJ2jkm4YVHAzSUYDrKkgnYbo8l7OqX2GkZIWMyVRKmNiP5s+JjlOvCUjJpDp21N9/f7ZGnIhQeWD
pL63RtEOuIHkMUeTSdpIvahinT8O/HRPLBAFt4nZ+/HsOMjy4+FePpoa1QFu2ullrrkdiD4HW9g5
xLhB+AoKLba7pMJc0WI4lliCnlhCb1cIATX80+xvt6grHhqRMoXyUe2bTQwp3F/0Tx1hvD9MuFam
59/sHpPm322/M1gdzPBhWWxDtm+HjAQoQhCkoANbzCPqqVv6Q0iebZbC4Dw+dCVrWdXh2UqMsl2w
qNc0dN+b/LiPc3qAnLAu6vKgp2jvF1uFNkKbbeasiPwFeuWm5+W4+HvuNxX4KlbJ/pT0ptIvIc13
1GNXRco73c/ISM9WAveWK7GMlhv9k6b0avM7FPOn9BK+o1usXfDgZaBgSiM6+Cs/49qIIQUODp6d
UNjfO9pDQuf6fOFZJ/7JPZiOEK+VvpVBk5E35XPtBGvK0vdIVRptEazuhJbYDcf/9MbU76mzlCyg
T+Har7TDpG0Mkr+3e2cA0q1FHTHZKacpBv5hI88sibaTO3RKT6QczD0pz5HTtGaLrKUJroWcjzjP
NBAGM5/LB7pjGkbtNqMWxuUOaQWQDDPgvk//JP2GfGK71AXZWiBUp1sB/6IYYUzcFgykKMwpsAke
3Y/+mURZYWJrOgPnpATwiExQwrHcjrf8QlafP01KObsjlLbM8jFXO4ppLdWw6B0/fWlKpPxy15KI
ZNoTsKyko0oTJ1AaL3DX+BveYyHoyEgzf31MB6tDwr0J1OVVIvJFfNja48ejgAPZyFdilpzPNcg2
FVLs7C9435oRbzVmf0SqQQGTN/eRz2IRR+s9LWbmRviSWRk6ytebgouZMd2Vede62DgitPsHbNmO
zVlgEaM1q5ZWP1W5tJw0XCa58+4foxhKiUHHIEyX4Y90yyYhpFHqpUZFKgVnC83Tc7/WmWmVAr/3
uM8+0pKo/CtB84460kzBNvmbtVPK/5yQ1P7kfDrVtsBfK8RbPDX8tXH8gfyvJn/KMrXPkRjudDzd
ojPcPv+KRBc+i6pz8nLbCBnqZju4BaaIYCsx7GDyiUEALL+J8e7aDXiVfvAYGCxUqgoWFUHX5iKd
vOVdrSxMrigHC7G0FWRRpCQWffYjvlmNkYftolr6ZMZCVtWSAZcVSWDjZKyZOWag0Ff2BTJQbcqR
tuOiKojYlG/gDPXqastvtAsyqGN5B1AFpaeb9WlWGEi5VzWZEVMx5uGvqF85YQpiR5Dqhi6nwk8g
KLYI2U8ZF4dzoBAY9SdpU4mLP3pJTnViWfwu8f1IYDNRvUprAtgkV17v6z7TnLb+7YbTyhIX0hI4
DRtfkWnUQN7L71YueE8OHaZDMY1Y0Uoo7D7pYQpHtitGfJC7kp7YihhyWIvRQu+Xg3syMGTgu3Xf
y+ggtRcv8ZH3EAPjXiEwWv/jQux5/7zKqmrvaSwmN2o074wVhq2Dk5Hj1KP+k+c9lv3R2QMEsGSn
KChoNYWNeZivRZsVVCAolWmmuwmwBKDrkN7OU/e9gakqsEmkuMKSDfbQC+XnY9DJptjTvYdkk1rv
8idlc11TzcJUvwsOfs0JjyQp5xMZLVdX8TOdwMf3m5HPvL6R2kbrUG/BaFN4WYS/Pd6RkEqnI1JX
1ciblzZRONDwi/sCfUVg9KWoemcKzVF+bUneguGfPd29rdDVMuAuw0mtDIQr53MBTG/UkdDYWg6a
LFzsPOjrxNokg2RzRoH0yHHFGn9KIAyu+WKAcCPPOwbs1vM7kuVXjrYYTLlTatmP8aoQ8TZQMPhh
fSAQ1bIhbR2IiTYexrq4Jq+Qi31A4xmnPm8VfQTAga9c4rQHFcPdXyGg+ITQE5ssh/SQ0mOZP4vJ
bkmxDEeqhwhUFihYhZxynu0HF8O/g01NJUqRcsKMkhd7q96g74dGZsk9P2fgbRlJDGfXXqE68TKp
x9TEjAr2WXIYcy/iCtTbzuNIJld+fn1gQqU1ekbImufhzMbM9cHgZwXZ3QuY5DfDKkkxtqaBqXs3
QvBt2tEfyTUKw/9jdgLm1Z1KJSOL+i5tj+NrEzceTMXlC2+Cvb3yZjNeuTGaZw0fupLO3LNP4ZRe
0GgWjZ8/RExTQVfn3dq0Zi4HqDiYZ3ZYhHjmNzaWJTGESsMAY+1NEhRI+mN3Ca7m8QhmV2GCjlHB
iMWlFC2SCn9cU91f8Hzv8tCSlw9EK3zTq03imZz7PWNEuuzw8sYoVET9UeucWZwdagVOHHT00SxF
ysxb9/iYVMg8tt9Prj/j1qZheEjySTJ4BujTSnUHCpYv1vRQozbBBCq7Fg3lHKjERzsYPYx6V6TI
U/gcLSQrGiFTuoqdkTTW/aFCLW6CpcYxDr+LGpz1CW9sUqwcijBUeq/DI2E3YYr2iH2/6xCuP5sz
XdjruWd7EqmG9QxRQZX7mm9/X6Bsxh9Z/7w20kM5kyFSBY1TYONP8mJz4p2SDqOx+cYgJu/WXJkn
SUBRv/3Lo/qQnLc7dzQXKLVmKjNlhJoDovbGs9Syd4eBzkE9DFaDbgVHePTusLpMzZxW+dF+XMSG
b5ZB47sB6w3JV8Z8/xhRh8xQYUIseKIUUabnm3QZOEPVTGqsuJu9Xg5f07NI8dTJgMelkf0Ai81I
30NDoPMVhaJVUo4DyQUj6nd8sbs+1EVL6FCBzKSxY6juqFo8cAXr9q9J5/LB8CiGax4r6wRXViZW
/1hpnFozRNOjQmRxVBuGXNO18cSKA8NIiG4tSpBjV7xXwMJzUZjoqGJVqah+l0urhIca9Gntdxb8
W+jAdWdzOHe20THtxdekwwoAxcSAcBVAS9ptzHlFlnnfJR9i80JSJabimgIp1+QpPA2ByouVzlGS
btZ5iH/f+zoqHlquwB7Ic5z4eiwk8uDygUJrnG07XGLxdnrV0SM2TeFY1DFvQpxMkALmfiN/pIHT
BHcbLXr+KQZT+E8+mv0VEzJ+hnc6thnhfV71eAHP33Wyi3fmqy6tTxmsdWQZgxSHkQ6bb5Utq/7x
NJHivpsxWmQlW8neHZVGSfmdKy4xt1mR+nUnrvyMdXM5yvEirYNC4RynM0Q2016Kt1s/9dcOnj9l
80RK6voobiyAArhoP5KPwTCTHFZ90wNpUNbRwgh2UkQCCQvR0B5RSSgmt7wR6s/vSfDjRoYVscP+
dT3q7SfHTe3S+yG58Nk5Xr+S4HlDN9mehdMITZB1jFJfFl9UeNpMkrxk6ija2LXzeX2UwEfc6mWX
N4sobjQc6FsaBZfQQqHKY5bC6RADmmDbrHIT+jezkLElL6wpyi6lk/cuDBig3ansE83He8pCIxg+
EJgu04DCMfAaRwP3h7WSVi587qOihoj7qtfZ9mPAQL+VjY/QiDxaTIm6Evdrtt+SN8v2PQEwNYgT
s9KfqVh5Bcp32astrb/b4HsDWNyV9T8qlKsEPuVBUpr7epSMqjrmTy8dpyAB8Livh1gsd88ocnj6
ZzPo3kgk/E+umyQ3ANfYGcJ+4wLXojBBpJonElp8FXb8ZvQAKr0BKHKdmrzYnBSODbB+zB79m+nd
s8EfMOmzqV36yXD6QJ372nLdMZXh9U+mWJAyfj5eGJ/oTksNTdauh0oIBGznSGzSh8Etnu3s/8zp
BXoQwbPGFtvAsES2POZLr/C3CZCMgDRYyHnaep7jWeMnHnO2S8KX935/61UtqaiON/U3lkQazLOg
eX0KN84SMKfG704DmMaiNMLMnWAulLXDQ3pXbKVH9IsVqpvtEaos4h7Js61J6h2dePcgIoXgi0rC
xF0ShVpnFw1fw8OJGMxITNWMHQaegqmZuKr+KbtuqyNPk0aGBlZ42inzFtbv4G+6pxVuRHFsK+qF
5W5UULMP2PDvrxc9+cAbqjJiiOYCijLWZ95IdR39rYhYaT+ny3KbomB0knXSf/VDlcQFjndxE67Z
YjFeC9mPebi6V8UKJTlc2zGhMv9tA7S4JhyQiWUQATL505DcKJ/tg8Kfu9x+laJguzrPH/rf865M
WuRnbB4qj3FeIM/mV6yVbHZTmWd5wygyAQwtYszauaERJ8glP7dR7AidpOYVFqUvJc3Lm4ocOIRS
b71zFQJ9dKnE3Z0obdj321buA3P2NkKh4MefrC35/01ZWXZv+kW5Q/BxFkA3B0GoQ2mZkWN080md
W4fPZOqMuUHsI7V5U6nyzJbVXceyMnSJyK5uPGsegYJCHELF1p07qC2zvJMQxvHdBQO6c+PyLrUl
9y+USuEPUFMsX97XJUym1xhZxDPz4VUGAjVffVTLCSl0npajV6KleRFkKXVQlRoE9o9LlcTEVtoD
bPKT5lO/AW0H83n6wqpe7OXMm35IXBWS1M0MCi+PI8rMzKPbTBsfXQ/uWvPN3fjjN1VtUuod1kOi
AMyO+DXUDTb1kgdmWNU05IShwr/GJKDyhwA3v/fEZ2XNzWFvoREMGYs5wO2scisnLa60lRgM27HW
Nbd0q8YQx8mDKUl11wZacL+VfuTmYY/K6wddzFup9sBjHImQBU9L9ZQAAmWcRKJuqtAGW46QiuS6
VSJGQjf58ljtVkECngT6zRZVviDWnAJh9r48IhsVEdh4CyGFpdYYP6YxLYk/+nRl1doflWWsZFM+
e1+UmnZ+E/0aKNl9n+e0tV0RbdEhAB6fTRhh5HkQRiyzluQXREkDfJFErpSyrsuUd8A7GA0j2O0B
Kfp9v/CYcGJISdM+1Phz2tW6/5heczV4guQ5GPHfHxFWpIkktKsad76mXRO5soC74qDvvZjWX2oz
nedJuqMwrITGiuNe5pIPwX9aFlx9d5x4VURHYx5lk8H7kwO3e8HA+svEYiVsPegYEpcUYuwW4mvZ
1sRui732GVbv5fPPftaEfj27WPM9pc21yETlv1yi98u2y6iM4rQRHTg7msI2CAPMoLEJKR4APrFk
FJL0spMpkK74K+wv2JY6tAS4j5mjZHzrG+3zKaRFunEjBfJKIDKYrdo1wHsmG2YUI2nrhR6O28ss
5bzUTbmbHnuD6Hm3oM+nwdTpQLk6S8Xs4+P59lcs6hMe1gUYSlMxR0tC5JR3NgrORy/sBLsGAeGq
fhz6Z7fE4HUa4xd2AYMoJyGzhT467uUAOWNtsYNzfIuCHERUc1GThYkAW96JvYY8TeTlYSwJpTZG
8srfJbp+sgz0E40UEyFsIbqGufM6RGSVEh+8zGlhSfQHfXung1XhjlnpEU5V4t3DPnZmUNu6YiHf
yljKBvZ1/x8hw9TbmoXmonzuc4phhKl1mmPTXdQSU3p2srkTad5JDJ5/F4EWP5fp+oeExRaNXhyp
Qv6qXQJhzPQ+a114Txij3BBGXJP5BnWWXjwJEjkpo+Ban1R5mI0a2+gyvOUlTOqkL/sbNsTVbmh/
diH/fiCw22Ehaw5uHxfWAGaKcZg5pSPSC95XAGT6OnFYB9j0C6HtwQDRMs2dRZrjYEfrfVxKjzJn
bZ3wTLTiOX0LCzbYDeRF/8rhbBE+oJYXMgxL3oA30PPUFwtooC88YZ1S6S4NQq7Hr8Ty1VgZHp2u
5vrfppmjQDSEsy66YbV7jZ8W+7m2qVy3yD1LIDVx79OMENCPRMk4TI6kJRBv0bcVRHHjy5FqnSZP
ufDppT9d28MmLORxLDk/lLoWoKlg+BVn47EDizYeQqktJVDfPW7b2W+9S2VZfvduzBBxqWhT1PLr
Scxd67i2gGCSSnpStGX4G4AMAD4q/yhQScWw4Qp47f8ChwCfsXDKX/MBmxg0hptaX122dSg8Prn6
+kdWSZszqODZsWjHxGWixC9Y/5gJBpHy6TghlzV6LMjsAnEy0CfdsALXjiEvB8jeCa+FOXaFfsM8
3sFf8N7NtwwZZcebf8SLSizvU26HWvawNNvnmfOxu+p6JgBDzGB8fiE4Nsbb9quTwcGdguA2B4VV
wBVb3PUK8JrZvxedyasawP+lW0x3splAFNN8Sm1bFPYmnr2tH4F++5eZdzhOUVb/5rTlw+sAJyM6
YAw1xStM0Zy2EFyq5OjhZP8UZAIAckFVKsb4MKjYdtWXK9VknkWXy+A5KfmZQg+kFc6+/Q5UkCQr
jfU4nwg1i/WHwZrjjlsKACFzgoyl4qDBNrmwI+O/x+mTeQnJy5gXXe1zJV0vtluq7bvyN8jtPPmX
6GwASkhta1a1NlChwpU6zj3QzhUQqiiKlWF1vOuSTRFTO2owTuTJef8jxZGahv5Y1a6/mlym+yNf
VsvKunt+I38yi7cv8pljcxohwu/MPE9th/eBQWaQsdnERJ9gTbRi4DrOFn3ZjddRTgY9eX41jUm1
+TkSk98it3qMMXF6kTJdbSEXl1rPLZrJ0KirNIen+GIc4hI9MhC7iRoYqGTIRbVCp5tpJcE7P1Up
QxxX5Xr7Y8ixFaMDiaTLenxD+WJxzRQwXdJAavSrJhwPr03IumG7CJvDVsyyTfeywOAQHi4Xt8v4
ZL+Gs4qvygZ/FZv3jIEjYG3M6G0NS6Tw6G/XzVYI9eGU66l1RnH4+G7zrps77QFTq4qaOKv+DUkV
qlqS7cX1vljmiGCfGKI0yfSn1ooftC5yY4bw+oenHfc0QvysSNJMSeHC+FV+M/lveMQ+j5DbzJKB
NX9ZGySOXMHfgaWdLNjSTyrcwU67PCfMhRa9a7fX96H1tj3eFzi8foBHvtnOYpnmx59+yLGQdQGv
vciXx0EjDDq1qFRDEbdgbzHISHD7Z+OSjZspFGnMR7PgMaBtW29Ukr0emaZR+stTy6eW6L4p4cn6
TlX4uCZply4C44JdoifHzAEt8cTnYncdkDSQiZmnnKN0Ys+G04i+msoE63TBvGah58wd9wXIAsz4
bKzN1aMm5jobvpZ5vCo6OZVp3TgrDP3hkf7IOIdeEnGGgxM06mjsUPCluv2yUfMRm2a5Hi0CU4Cr
D64qrQOO8cODmaEGKDu6h0zQHCTouQXtCydRgN82k7Vsv5166Xk0isKjXVKR6G6LsTcdAtMI+Djo
biLOntTA4DWMOKknUgXAxUx5JF+I5xvvjQP6UFyVRXDuFdmerjT4GLoftBvD/xEUct5IGzU+Quxt
w6eNEAy+XzGRhKUexNHoTRgnM5cWymHuVb7izoNFv2e0AZ8lJd4EbGmLlwvCdimbWXPHkb6HT2/2
hKR/Pn2vTAcQ5kbR9aDgoz1G0RA402ggGyY2JD2gLFrp206zFCiiy0BzEn9iaSTi6uRw1YtnVio5
t5tr+2mrDnzoFIKlzF4lZC+3lu/WsQouHIVbjC3WvBI7lWmktPaSNp1PANQXOkqNBm0Z5bEp0Ry8
J1nQXaJg9QvmkEC6kmiXXjO2nORYHzHJxbJew5x/NFvVx5q3Ao8wkB0RkfuhgtGhaCzFlxSeScoR
Xc5PznI1hfU8Js8GcNK/Y7sxznW2zJrgssTYLH3ROcYXFmsBNU7P3Ygu05zBzwG9McKD1rFt52oQ
+ntDMfwKyJnLXT+AGTEl1G8N82gZwYulA4zPYzyp3putzLnGobHC3GUQT6EVcYBCFL9cjaTFzM0G
lZixjht5GKg5f84KBzw7p6FRiDKPbwkaKhMOSjHzhoExFtOULsyLABbvbolN4gMkBybwmjRhwuOU
LP4CBEQWTolaEsWygprySjSwSo2c444nvIpqZYhJAn/UjLpug0tezAD4T2YHrZsfGxmGBrz170M2
iIBg5OfccP31IQG4dn0UVNZz6xDTIrPB77GXCobjrW6dP9gtGoR4m7k6IIPpcMcJ5TL4tRKeSWVb
4jphQ9iWZCZA6Shh8dG88qBJgPX+cPn9wlsgjfLpmn5QM99XmHJQhFTVhN2FTOIGI6HsHr3myl5x
xZwv0WftiOVGOvnO0CHrYGlJflzVgavQeYb2+EAcirt3jEsndupXwtFFGeEIOgPzxCyl4tgAl+a6
te4tgAP/+nFdk2Pe/Y40Zw/9xsyA3/LU3JO+8MSus/vULIghh+u7cjDRRsr3/fVQ1hYa4gRVUT6T
sePq+tkBaGNxb++19uF9vVMTzlJfrSMzPsYjQL8KhNnKOJSijHFMsoHDvxij/ieP/YvJ+l+q285i
QTJV0B5Y0NppOAV9Z64jlfJiDfJvd0GFuUAmcCHA5R/1mXHPBm5ZxOfT0ZXmiF2E1zoTEGQAdtpR
Vx87tsXO5tUbE4KgrpE+5JBtNwpLhpwORxbjOHtul1dm9f/mhtH49gAcJpsZ1gwJG0oAUV8Rzagj
p33gCS2RbNEghIEa3wDqSnT2ZsSS3xzWPQFuzWlNs2uff0A+XeLBBOt94HYpL29Q5InxGx5A61hm
rhn6fcLLxXv0zevbqd4lWItsTO+PpS6W7ONlCvv1TB9lDG78iCqLwj8SFdmKauhYnIw96f3sM3sK
sD4oQdInvs512/o0VWuUeVuzP5HKV0RxoD+UJtYaSvvh8WFkIPNjZgjdxUXxnq6MZtI1K2yXEx8/
suSkxjFdSwg4wCJ95w3wzvbi2BqvbgD+rH54qqEcnn/3OpvOuMtqvLqxCMtyMLR09rJq/HH9eG8v
JBMsnhL1RHF2vRGPGE2Ewhde3Q3UxfhdfJz48FU6O2iibPlzlI4xXCTASeP1ztUouCy+glAkHWHK
U4uDmRBtR6c99yZcbckxtfPtRx9voYpQDzstroh/oYRO1OY3pd91dBcSdhSJasxUwIc1+jD7pEc4
UiDchhqLEdDoGHhP7kkKk/RJ2/r0NT9k7zjui4n7L2JFyb2DNE/Ba5g0qYA7cGd/uzQT1jPMCnv7
hbFpq74X5SBxqtCCiXJKSpzHe5znIRvEPnXdVxdnVQ0ZeO2+pcAWxZSCuuH3JbPxX9kbRcByUExU
rptusEcPLh4rnlXAD0BkpEoSiEfiFH9/ZqT5NuUzyrR3n4sTIDtseciPxF8j9VLJ8qdpkyy2U4h6
CyQ0JscrObYvWj818Qmfrdya8lyoDd9ujx/VwoD70DUxTymBB23sqhSJeE8bvTPkmBqDQ3Vx1iLH
G9OEWJ34EeotqKBdfp4GeyZ3/WXCTA0wnge5jPNbG3hrggn8cdMLbt6PZixEGQkwIG8Fb3FKwqps
eBk6/yg67+9QNobGe7JYJhXz648AWye2os4uJThEhI3tBCodApuGeg32s70ExNur/FKe7EA74aMm
BR4uWGFUb4i065T6G5ZkpaYy62xOPHFQW//dn0OSyrLk+/aBxXHQu/KYz3Dnxk+KxzNrMo+ej8Sq
UL1plvaZBekEPEA/DGYi+vrcS0Xg04k3SX5T9lYR7G3xcUf5txgbQgLSRm8OoUUuyTTBRDJrBPuX
kPOrQRKR3pm9mlsrQ28Y2Mj+oQYCjtTlNCChXKYCXlmhGphIh0u5ULharCZKO1MUp7x0raDeUyfI
qTr52qBwaS3emiCXC1E/fnaHZ024exQPLDxXcQpiR1hscFkLeeZ+q2bVw1AFrlbwUOoKuk9WYnjG
KaXAIXaajvyEAq3cD1AOfynB7hppwI2BPg2niYXUhiB+JhdU9M6cbSfY1s+7AqIyrIB0tlSXvnU8
Bo5v+MqjK+NEv+TzEWX8EmDYmtYcA/KGNxiaMCBcNQCjAbSbBAt70V9Ofukjult/GSB/vVSRJpVm
BMSOAi2R2MufxiahsSwG0AqC/bLIvow3Rd8VvNYMkNZ9iJP9BWrjTj1lrB5FmS5mJgMmBMuruAXh
BM6/WMY2dO2mYnEEzRzVTyjYFckG/vozVQRlJ9uqnDve8DjPDI4Kw6jxJ9jFCAXZcWCvVmxAgpzz
VT8xEkUZPMScTdE/AW/EQ4vDdf0PD3BFCKaAPC/IR2HDCfPEGiuZ7+L9A2k/8a7j65Yu5L7zT4/n
MHpcc2CepkMP0V+B363ohgew1lDW9dLnNsvrX4J5oCLA4AHPbepKRqZCBrjpqcULzXAaBA+zegVW
ryr4BnceGYlTb8N/kJEV+6b2487h9VLGU+cWstBCuPLXQEOSqxS6q1VC5CtJ4OhNu4md2TWGE0EC
lL616dr2oMZUoNh02OPTAD1mRAabwZipZ6Oq8pW2AEFOnEFU1CKxue78jOp3iR/tdEqZDtQpCO7s
67G86sI5aTu1crlXaY2c5ToH4/JNQdlIa8H1HB1UpScMzm+07kbOqyMcohyHj2XrOyjmQWT0E6bh
qfui5D6DE/hfi1Cqh8eOOhBYouLQhou+gXnqQUrhj3QJ1+h85Qoq5r0M9bYXq8gfgB7KaVWcxZak
CtW2c+0+dykQgAej0VF3PDnA0ukqi7Palssh7CgCMp5TP6lmRLFvTxl3t24iYRN/JrMC4T1ZNAn0
+LFebmcmUD9Qdo0cUSkF7cMa2cWOx/seGpw/1xyfxEYUc6/R1kkkEuhdlS5Uvnb8vSJ4kxfy5TPp
F8sWqoXAsE6caTCRnn05n9ufrDeKMNLW17aO2jdWZMkyCfpwn65y572sViitVIHwlJhuhMEXu0t1
F1MXmOWMAclwu0ilVax1Jfku2jLYq2abq1Bhl8DxPKWs+NaD2PiQLD+a6i+8dZaJ2kTXrJsfLfWM
LIFeYCHTqThdZWZte8M8VyFEfzwDa4tTC/gYovjEi8gCCjg4ozGqpVqPJWVGmlYXbMwGNYeKMqtS
CGkcE1AxaRa/jP3Boe9UIY46FWY7Zr7xIsoJ1n7Qdr8BTKWAqDjD27O4zelLb0pBGSYq424/qGT5
+KTUA8a+EvY8npOS8KtvU/+vDBggGH96soAUVPJrYG1xX0pLOfACFd7CRDNnlh72+NPspTr0zpqt
uDEYgs5U2/gMPKSZILBm7pPKK/sI1hAZupLBGjGpNyoPHl1P9CM/4wTj+iItLc3af9uiSnnIPcP5
/pP20tx+DGwakmPD25kIF8eIsUcegYSoQonuc7lc8BFwQjO+WGqA9q1wsJ/RTrKdfznzc6FLwY/B
u0XFIJr0ndiAbRmutDJHKUrM8pNloLmL6HICm56MM/6zocRX8ZzJ/7jpdzzK29xqW4DmmBAHgMIS
tFkQ2PsIqu2inxaGsFe8OXbTeUe9QWn0j7gao3BwwXiYgQ4nO3vt3Z49B6p5Q/aOYn4/OXKvVKFG
5Tq6d7VgrDxtFRq6jvztUh+LjcJpciorll7SNFS1W44CrRWSuIZ0pdt8S9vT9/Dbr+MMEJr4m4e3
t146t8ulFsytZNgHogLIpIxm8p+ZDl1UCEcOvRPD8ajxXfTKFBhJvzstYjQowmJHpqLmRcNRTwCE
R4Kp3JQNNHeM62JUaPsHA3b0/+bixWcu8YS1xzRhenRsEFq2JJzcFRnlzLphgBgZbqhi86zIxQJ7
SEV/e9/6RfxzkxcekQPDTUZw5QBssoGJnAXeaOvbj+wNEOuTK0+L5zahTnxYPeqnozt+oNntk25Y
dEAZki/Hqp4VvR3URLHaCWUALx5XihE8M2Tp1ei6A9cYTH9bqmw3VIXcF6Z0Xf1j9LOa3EiSYJqS
XJn7JNp0NaSTrBnf2R3OePByqjxmL6yJ5TduJbgBsdGscN01ynDGcQZ5CIlDXoB0BV42dElV1C2k
n5nTKG/h1mpyttu/Rqhk4t9kqPLXhUt5K1xkST75v9XyJxqGGA6XDUBGrKSAK/9Hjdd5vVLc8k1k
ujTkmnxCCKjxYXIXI9pCrqzLllN8eoMw4gmvA2rn4Qjr97zTi5SsqO/RBKf2g1lR69hb22nOnh3J
k3qvNXa7JTSz5lZnWbTEaFCMPOJhHRwJckROGFfLFmUES+a8Ni8G9ua0CgG7WDsrDM9Ym+YAYdx/
OpdATnDqmwYaL+bpqvbid7jsGaQzngvZlgbXZKgzU4UQWFT9rNh0GW1UFiWfbw60hMV8uVeYWvSr
nr5cE6c7VJssPqOkZs2UDTkBtGduFVIP9f4DIYYdI2DB3nZO1hwh3NLFKWrBhOSZ8D2urwLH+5Dy
3G/7UHtk+ekL8iLLbw64R04KJiJe7hoOjzpl8ovZ6hE0KM05c4RpZEi8IVIb3FebZnqs175P1f7W
X5mdoqdLjghIUrawbzLAEdt26FBiZXiMXKXz7twhUJw+5bR1zHloCtPRxXXyqI/brNkYKicOofBT
FIJZO9zAbiiip6ep3I/YVaacHuUw4G0GwbshdgX8us7+mxALZ1oGAZKDTqBW9JwOjNcux/t/PVuH
PKEHZVRM0CRUP20g8GHYLRIczN5yWT9Y6HBS8evb2YHGgsAs3ZuaEP910irwAo7SN7lke68KZ1FE
HhvbG2UkUxqXiDbjWHJIpav2zVlJtAOrnhOrRxHTE/GlJZn097tOpezLY+HwVDdtsQ7BHrv6GjEc
Q9/NB2BZh4ujVfz/WXRa7A3OQmsRgDi72OLrofvOCxw0mCRINDvsclq6kIkCK2rzFNiAE/DYjQYm
YnxyZDhya0VQuyh0LG3Ei0+dQSfMEPSYtWUEpUNJY4nFqImLz1WDNCUp6zKqKQNLDWWWa/Fel4FO
A7MVNwroi9obfdICIDbFu4/llHoB6ZdbEGxYxIobhXhCXTd/cLAB55GQG5Lg9JddAQ6V51eYTYet
Muct1kg4NiEWEo3gH5Uuh+PEvPwLSvDlFtOuJQ06KfKxTcSvhoxtjbG5981EArFRQ9+EIfTrxxj9
S7PTxAPupFrzucMyssUhnAQUewYmXOz8k6eE8kj+ncofsatSzD5Ks3W5oSY/Ifpex6NFrggbpzHu
62GQTvN/Fq6xfegvxqM4RvE8boFvrgBl8EKdpzf/IaQDZjT90GU8Oml/UtbcauLJWz/zsAEFFFLs
VKB8WWTvoscgcNdF13wNhEqEf+JykXdrD37sWv7Nu+7IuXOQn8NvWnSDmMkrsFqOZ3gKV9Wayrsp
zFeLzm3iElPkAwuNeoN8kbX8YxZFcrE/v8sSe4skf/7UljFn70UUARFrdngw3GNLKfbeDXjrR+5N
QLinkgkZcegEg54QWMQyoV0zcr0Bg55G5q/R3bd5QqFYa95ruO2VKP7uBE7TIOGR4phn/oH18siI
8/iohwIVknEyAH10U1a5wCc/dyQllRzp+12bBKECEpUhV49LEyfwWxC7SxwX07I9Fio1LEhL5d1n
ENzj9/BuIn+7mWc0PG0/LYRwXIwgll+GFFoW7hqEUC5OVI+mdkqwnh+T/bRsy98l2FsIsXfhv95z
L053NKWDZCHk+VgIosj//9PqdcAVxiLx53hf4zopnOv4FmU/fGU9zec1J/J36rbBhVt/iim+BJ69
CEMvsPW6Qj3UzjNBQLZWfSYTRa/0YszcewpCT+CQF45Cw554Imdc5QNmgET72zNeqtg4udNby/t1
3LuQsPB64hZAm4EsfmagPL0N0MGoGjdjJE6oirfWDwqw5UxJuXtoex9JCujv67DMI+3YBaH6wEQk
XanegETNnFkARkV9ykj9IlZWSrdA5T0sT6HeZGwr3pOO14WNSy03zpXp3OREMC0zFJxp4HhTcf3N
mUGKl3mnx+yd9qFnz3xuDc4Phe8FTPf+5dn6/uJksWGhuw4OWJGQPs7knJCaoTzYIP+1aZcX0y81
IRmqwuwsu/XeY5DcwkYjL1gU4AdATi4dpvv/6ONEDpPFtW3LctoOinBcIaQ/+Y8ngnNTpL9tzNIe
DWJDmddlYOQZr53ph9PZoUmgsv3xKAnDZwlVxYfE7G7IoydutNUHEgBXRH3OiJUbLUbs+6nyC/kM
7a11Qa4osRLFEQewoO+zOvYxWOlBwYdtZfzXagZ2zhllGN5iVQjJ4BPhqBz5RrSUKUBrUkUy2E/d
RH0YtZ4CPy3OF+bc4jkCz41cOpzsqEAlzw0p8t21zB4PgEQh9M8D+Zjl2gbXIrOrlQ96CB5YNoG+
drAZd4qN6xE+d1P2kizKo0dMVt8VMLvkA3GYoqDml+oPLl5OWgBw27xLPrDc7YyjYGtkGpVGvPRm
BgbIwdyynDyproIkdU4z7Q5lJJJrTRnCKxKhGMuRuJUhqTzShQ2pS6v29saIanC9BFVOWXFesuUj
u/fXULyxQ0VF1vjSxZ8soAr0CLszHz4rZMbrrIbZbKQIS3pEIZ5meQM0aPctQ37pp8vrJ6rgVW87
4I1OqC7f/ftCGwiWv1G/WOeSFCnBFQu56qvRm3/HMwd2pRBI5c1G/pzeDrVkTGdiSbrOdEJtB/si
q1GyuOSTnwEchm5lWcY3XkgO/ANSGxnReFEyQDDa/P3LF6QLcKOMJfkE10n5n7/pJp2noWyzYPM8
I+NDvmeUsSh3ix6mDj9HbrxABaqk4SuJ7FO5tOIXLgrSFWCOXw9VzL2wydNZUa5pbPTLz8EFfnrn
q7yTRPlehHhrI+HvpUJL/lw5XLzow8UZBi9gHp4Mke0gl+qpxWYt2Ti2A92Hpfo4fTOV5A2qTLZQ
ok3QN9EsBiZqt6RbIQkUbOFvPtIsFWI44iGf1ne3bPcULX9PwQvXbFGwkojn+5/2+Mv89NtSJzo/
3dT+KMeStTrwAREti0HjttD9ksEFkY8BoPbumSrPKRwl8iHvU7TJ3OyW9K4aKHVaXhE7rYnREoHL
syvR1OWUsW7hpdwJ7kbtcCZwnGj3DHinRSgyGcRZs+BkFYI//g1nVargEax6wJDKqdVcMIFW7mWM
1s/VrBjbMtbJAyT2qmN7AWRvolCtYzybRsRkaiYSnzRlA1xNrGVDoHcwHhBPe8rI803QUwS8M7SN
6FmOuAVl6zG2iRS+xXswzPP5z0jMRNO+3iDjb19iCtJsUFPVKAZD0GrJg9kj78JTTXGbxxibSgb4
uyPd1wu72hefTljL6u+FTeTiIwEb9BoNI7ua4d7Yp2znLnRBpTG8gb4qjz/JVcAuWmmPB1gMOmIS
egeEDSekNjoR8RhZu/fxS2qU5B+VAOJ5Oc7qeIb4pF7JUPin+fguAqYtzYGJlYRt4v7APAJT++i/
uRUm0Ju9OYy0WVrN7JF4yPP7zz6Cd+yq6FnPQE+HlLLmTqUqpVacSkqpS6yHu6K/S2CN7+kBbaAM
Py02gaQgprhkGsSVEhdePRCcS6fzu7RNDlC7pitoaM71SK/GYVODh8aCgBGWkrRhvIE8YO7rE86L
SpmcnDQ7hud5sKpNkqTt4I4DRUI1GfojcMy8QbdqGwjNDr6XpHhitlvPmAuZ+Exv/7Nrs4E1xINP
t7AsG0wPztDAYP0NHZCHsIZvGyHQWL5uTZhOvWP76agWLvWIfXEFFyXkrA+h+YI4CN1QsihydsHZ
0tiQxY/i3Ch/ynZMFJxEcgioS0irgLmiMuNcMo8LBFQpcsEfH2qPUhXBvoQvoX4gg0b5LtuH0T9q
ne2BFau6EZIDss8aOS8sd/aR9KGhafJbvC9WPbIcpDdKBSypd3X8SVFKxoLde7S86Eju1Dh6Vl+Y
n6UtWyfbY9iZMunB77A+IXcPVKPCEpLpQdj+TKexpNY9tuO0PfhUNBewgnPkDrYWCyVgARAZirR2
sTGir8rriitDH8MKPmYhv3OTsnaInDVGV2scvIWeKyQGbDf5Dk8a9kmOAMh+mnPbxXoglvWS0Xyw
29210IOMxaGlRNOjJeWXeav51bZs0oxyzNlEgc9UGTjgco4jLgl+vHLR6zswwdXi4TW4HGOqpq/O
pMVoO2iUJ1bXRtYNhRjCS2KMSwjkQ41HYlM4/uIGlt0wu5aDqx+GE+h+OovV6hufygxBOcsRmQIb
V/BIhNVOotUgC4/H/0D+YsxxxwG92avUCDBJiYzVfjEcfI/WnSTl4ZHCJ+IDrgCri3cvnWcTbf3b
FoU+OGd+xA9Ucm79iHBRgaderWq6C9hHZTgRY29sRWHtp9leXsmLWXF2ynJ4epQSANtZk8s9ogYo
QRNXLn3mgkB92kHn/vLZaKfPdHUopnG2tcGWkG7x/sOafbQ73G5U4Tyzud5codjaR2Fwt3ajdoEM
1reYOZMDy15794re4RPatMorbx4g4x3JPHv0QuWk2phfx/+5Q4/QiWhC9GAMH3IsAKsxR82ZEqyB
deBD7NDx1n/kKd7a5p7FS0x9AEH0P3qQ8HddgIpJ/Gopri3tmTRms5n+juo+KP4Ik+NgqUJqXox+
WNt/TLM+UkqZmKDp3Ow73ScHg4fh2gSl1I6/gze+BMCXNJd4j8bvtoQweUi7hbHcwt3osGyReVsH
aV7F0gwtniz9UBMRGUPfSIR8peoKWAIvhCAUVgZGPwARHkOrByKGG6+1tFDeq5O0HYQWJ83zgHGl
u/hiDyEYM/79Rv0hQarThi0QXsSheEdc8h4sd+ChN0Af4BKlRT6huGpnsKOz/R/pbUPeOOyIiWDY
k/GBOmAFgxJDAVjvCrJ4S5gIjKXpjxoAHXjVZ91wU+vSBWuV5oYxeYG1RWpH6lbZySVLIXhb6Xst
XjCZ+GDepSNJjKcsxTv+MDy4i6GAM1ml55CtO5ArcJobITuleuIcyIY+mxK7tTLAoXQMaNrhUTf+
wne1lcO4nwK5aq9gNV4Q4c9PTA6/Tkbeggo+/taE0uNaCy3D+GSBiqD9LkUeXuKcsvUEgw9NJM5s
v8XnA7CvDKtHLkBRUtVOz8dcPY1zSCecIAX+q4GqAtxZuRGgO2V2c22F+jQNWKYe1E8VlYilQbBt
1M67VwqT811aUdG5QVE9/xfuQqceD1LPuojR+/vNVTGlnJvgqF77/BEyXgYmP8aZhyAawE+ggL01
KwmP07hKPUWXYoSEdAgVV/rfXin5C1zJ3urLrj1E6GkNjxHCbuNsrsDaxmejByR5OVdn9SDyRXBe
vw9aDaLkVhdi2ty7B6j4Wgp8iBReNvljJdTR/1fkRXLymTr7j6/Fpta206oAgQiQLnLTqKG9l1Yi
2sqcg5PgjhxrUjko6QnHuhkZVpcy/wTrKcJk+nEY3nZ40kkGUH1/ixg/ATWSpUXtueLCugEKmkSW
INxmQuGP1cjrKf4LZ+6AGLP1HlsJ9tWuV/5u8ce87/zqML/8EjwyksYb/F+eT7ApF5xVr+Rih/T0
moWPrWcr+3j/mE3Ug8DR2PH6oa+GX5Cj1WN5N2fBwdsFHzGGxEEPL2IKSVCDf9gmy8QNi38iyyfY
06R9lHVjUjfB0UwBtjp4HDkFSmNKDzBQTkqbytYeAqvLzaw959c2EN/iV1BrdLPZIisAhSHxIKkt
WFoeKWfEi5oMv0eEcNEK23R7L8HSuByw9MATw60T8u6VwYGraAqPhguCqJyVIPcaUTvkjktCH+/m
ZkoZLKhgGaR0EZgf/qCVfelT9FC3GbKaqUZ0euvX4d5UmDfw9ND+exZsv+nvoEes3eKKw3/ovj9E
Ps4bRPtCOHC1JmYBps9XeTWDXpJG0yyvONL3vbE9dVUaDcCUV8/njIakLnEGd2f01UbIDKjBBtpH
waqedMc05XI3zMapfMliZKiH2Q25DC9Tre46oUmwF04Gm9MGxcCockLyOmkSyEC3mM9XCMcimOao
NAKeUb8/3984/rzbLaXO8pgnF5VAYbhSr6j4nZOHhOqo6vud6VWHwzZyGi3li1Xfv/sBy9OLDK8Y
9RbTV1+PZ4FRJ8KtaUk7lxcyA92hhfxUxYcisipJXF7y+7Xnptxc28EFEsWNovTL7OvsexgNMNA6
PgpSVtV21K5DIMbbtySN2DnJBsKpoz1QNPnCsUYq9kUS8C42iPKGQExEwcgIBD5/3vrkwmpFMbmI
58T2PBk4d0pSzM9dCASTj6yPYDNOjES0F7XTeCC1EDbMbOnMWgNqHrbyDXj6a8SoitnOI3DrGIPs
CikkN0vsTMlL9A2nfBU0cRFg+8yZwSD5QpmINMED6uXvQcWdmYHmuacGumiYIZo8DV7Dwx/WP/26
QMbcfN4OYX1UFHNnr7VYLmm2XImK6iDOT0Uvu7veqOjM/QTHq2/tymItkwesTbRLdCCHvUl+JXEW
AYDfRGJDgzvYqOofYzYJxVeOFidD2XIB8dVP64kQ/PJDZjhHXGAK19fzg9KhSOUX9IXGaRyzfzio
vJ1EmFDxOpGvhyEpPNNXqjIFo+gknHP9edTnZCX4xsVA5GRVykfaiX7gfP0wyJ9rM8+dKqYzfHp1
F2Sfzo67ok5e9N8u3fSqV2wLIUL7t6VFBbpgNjkQXzWYU2YkjrV7f/QpXrN15AYDxshALhNhv92X
d99yGRvj3HVtUGgK1tI8g0q6uxcFSGNnU7ASaZQBVlNVl1ukqVYGS1z9ltLmgSEViqe+ICAAbP37
mWg+EO+gRZLr9AwQ2isS7OwcgTSpxuLASSZWyPFYxpEV0h1+CS7Ln6fys3qj6ow8eB1GPoIn7T9U
A274SCwwYejTPT1r+0+Grh3xRZTXl35AjtpxJjj7l9sGX3OddqgIhwW3jWScWJ1bRpgJULbAq8Gq
Z3lPl1LnKj5eu+8p8NRFXOyiUkOxZfpfcLjG0BvJc6wJjjlgfOOGwX1s0Iq81Ix8/eEdsqXe4u/E
wV10hrQ/aZBRfWsB697bQN05UHHugjWJNloeqxKQzn3MKH1NjipfM42qwKPIbfhxDyqqPS18aV9v
nMEY+V4zbzdUp2eErvc0ymh2R+Jc3MTLXjlXrfXT3VHNwh9pC3ft8z1d9fBDGsL5L1e7NWtRYu+R
lspTPETi4adlvkTbdT9CQ1AxWEbw3C/6F0cEHZi7IzXYJ2VsVK8EPNIo6u7EGeI84EOUUQgvAZ7O
6O6vIY45zCeQ0M656MuF007MGYf47dQ1iQILAlR1rHBqPKcfmHfNXkAVlYoTFz5ntJOOFTqgpnrQ
UHYFnO0NF7JGWgyQaLWGgz0X79KFJZ8Y+RdpAP3oOVR3iqGCarNYYQvYzh1m5sdHgZqV6hi6KF0n
LPRTYwyDCcFYlx1foFAJhGrquSPcDRtH+UsCp5VxUiU4jQj/qSPn3q49gFXK4szBWKg2PuaT+ivn
0O0sdt3T79fMlwLdqXLycVZluORg/YmpFcU52RKQsNz3EHM2b+yh8h9CQXruEHS9FYS7NXZh0W8p
cnAoNFghoUzahfq6pHjnbQuYYNr+aQCmzadS1WIz5Wr1OATp1793iWvSVqmfMbM/XpA3cz/UUg6E
FOwipa5839ymxNxSuC/vlL3vQ3b293fZgswcwq5ENL6xREmZ4me9sPfCLgUrmYIz44CIisOB8CYd
JUp5K5tBxkHpfDen5MPxlTqzXDg30v/gflI8Hhz58lqbOSIQuQHCFfpnXar7ge6YIeiYhQN6I1fR
fcigjBBi63c13GQobTQD7NW2Db+V/R43ZCzeH+UbYgBhfgjuVrAV+5DCpmAGv4mbTrfCgIrbypR7
mW5Nd6Vask7jMjqL+5gq2QRR1m0C7N4NFCZj2qKNlwBmmHcE/N3NCZGqPZQ/w37afdQo1FiRerS4
4ntu92rUm7NYM5NLb9TiPYjoE527qf83ToHLEfzfWMiYYQ0SjW45zKFsk1l01FzTktksssPTjV72
7D6XZ0OnyvmcOVqDtRq7//jX/Jsw37/w1ppIbmyvkqs1QNNjge1h7q4YQK0ASTl6jBYcvqcD+dYm
mkf32UJISW+Rdbe9f4SK9p61HjokHXDBJjy5D48OLM5UdH/yWJzsYh3zl3L9ODjmAa78hNnJ5Xu8
07dotAsxgh4p/ink7l/TyOPeKIojJtbFStlOoD6UA2u4vB/56y8tg0t41mPdknnos6JtWBBODjw9
mR6O/+Lv3xx/7SlJ0l5SorKJkpwxGzQ3bIlwyD2mne+kLLC3XkA9fYitZLDQ5PmV328KBndDZ2sk
kZFaji27p4DN1cLEZfH11HvnWwDfxzqIAyvD9ibN9MTjiGO4AsnDkuW8UDKypyAsdbcJgWw8EWKD
9oK4uHeEmrDmowI0OkZ4pXw0elPEhhIk3muno2JZVixt7L/jh2Wb5YLP7wvil7jIrJdwHV+NzJtc
Tgm4UWnrA4QoobnMUMkUgLHHNuWYbN2ftQ9eN7sh7i0/oEPkzqtYGq4ef3+WJsdG0eiqxhNJXEcA
EFOjnSpxaelbeyjigT2bdEALUzajmhdgrdshknzY3Gj2gvXoq85n8qk3cG9CA54+YWePcxunAch7
V6QgI5T4nA4U9WorPS3KU+Ml+gpjcJwAKxU+7QIUHJpNaicaQAAcjzIwWVEg63TjKzUDR8h0z9RR
98eoQPgB0unGi8mVD7vu38XghJYGTOx6o1SGXs0BP5XFpC/waLsrjNxpBiki76Ummg3wO5NT7JtM
BcoRP0zGyBXaDIPtyrxsNrAtq21Cn2SjfW8ibZCP0E4unCn3h2O2goP3UGeZ/Umn8LGzQWDRIlg8
250ZEjN+MooNqJTQfXmHxXYq0UB/HDk84EYUD/n0mv1UrZEFebArPqGvkRRZ5KgvogjBLjTUUA66
IfymncugWer99OdegOgV+ToimEzX8DzEjPxlzYtcUJqNA39+9WT6W38msJEzjU6fLNEvDMenNC3r
BZOCW0jOJOP6prgcQKbKAXGRSacD9y9xzteQ3Rvu95/3Azq4/yzkD7SNtPMIT2L7nbTWbUfUEVNm
3A8j6xjSSxddXWtzebQak1CJ7OOnfF3nsZDulWHbhlbOrBHS5MGoN/XpNXKvMlfuvmYNRjswd0je
H2sG228U2I8fMiMgmDzTZLwZ3VkQ7JeBbu9WpyIO5uc+2Tp/oGifbgn7Wc494+snIbmYyf0Q/fcs
Qf4QG5RGrX8QoyDA6vNnXb4DDNXC/tlMdcZIX4Aoa6J4CF5gzqfybXdcrtME5NG+hcW9PqNKSZ4Q
JoHXNaSsdGYO0UQzFBAvo6ynyS4hHZXkoW0ctd2t01JcErgk5wVDkP/0Ki9vJHvtEt7GSfJ3xabK
60idKgzJIPffGaVSfc1b8Mc9GgbyAEOEfXpkhOST2KNn+vmpL9ReDnyMMRsVweXpXwzwT+tf1uUd
5RH0OPLREWglE08kj/vPkZWagoB2PkNGK3+Jy0AyVpEMJCg4WByQChLxkY1MSQhdSwPAb+ccbSqs
/FWB7u5OBZ68VYMturWwwVNTEY1Mx46OL0cCeHyGg7W7flTHj7DejdZ4o/3xYR8K5kdnyVo3YlVU
CgceFt00gSKIwfzOrWLzxZzUAEwYPa4FyX4NXDEolrkPc5zbVBUFgu5uF9u73yYg7lV2ExUlhPxd
rj/sMRd2QqjSooJScKksHoC8Y5KG2K1Pmai8IkPZw53BYoveexCzC7MmpWL0IMFEgzLlFOFfZ1/S
pHwZh5mD7o32/pld+tVwK/Styo2uFFaIEXnBD6mdw5R3M2uD1yHo3B6PzScAkVPZ2wdKVAg+oLbW
zFvHbMLUcVsWT09U7lXSiS1XM94iqef4xiWDq4fELXopwNYGk7HQcbD0IfjTs/jcmux/y5y+u4es
aLxu+9kYPxmEzsHjL3JglXc6Qz4NF1wzmhk9prsjO5vwxEec1CZ87Fn8dYMeNmvWxV5Da/iAjyXT
e4Uj6mqNmVP0bQ7xWC+YYtHIP6o9k4LUE+PpsmwjUUp3QcFZZ9N1XeyemucyZNeZCUvDltga79jE
s3B1hF8ihjHaUNuANMcbHHK9OxZgm+nZxlSvjSuHoaHn7+ChvzBC6ZE7g6d9nPZs7YM9LWgN16iE
AXqH5sfZmgSNbhMk4HyCF71oaUfpO9BtFpZaLlC+pR04PYa21iV+xqisN5ok+G8RCWOUoUWoNIOG
MYhWX2Hqnzk54wzoduGZ28AvousRb3nD4B5FsvrpKvVQSx/2YSn+zUX3ZImk9yMbkXl7z1K/6MoI
eaKLBqHCoam1uedNFgoGBGXz8uxFxedigULIAkfHy6tLwpffH8VawocQ0RxuMiypLtw4ry7942mT
3bn8R6t1Aq66fhz+vYfBJ/Za/fgJFgvdfduV9GRPV3mkiAOY0jJjfNHUT6Tnm0TBaGvA8RXYYAgH
L9Fepccz0FemNJbc4E1GM9HpvF3cKOO317cqfBtrMjgOwzWhxLtbHd02I7ksxVnj+op2MGoMoV2G
z0c2NC4KJgV55C3lxuqg1lFRVa0/9zx11JIAwLx8Et+ZY7LCeNLpQJ9hE9FlevLBYFU/flr+EaYM
CHJhyL4ZR0Jy51JykJ0at0n3+YODAcpBk7lzts/GNqmLmjzyuKQoaN9c6rzoUiWaQ3JAOv2JzrQx
NAthiV176BRfEcHTG8IWYKjnTkUDImMNbfuBQhQx+GM1c9ot/PF1bbELKAVEXgaLO5zUpykpMNOO
aUO5DVLyiF+sE+dIqMqE67THrVaslxCuRWTOxb2Ei6YMn05jP7/3hnnJA9IR4aWh12rgEnSrrwh6
9LgjkztsxOmor3Kq/okY7Iw9ku8TdMZ/cMEZV4xul9FiI3pqKlTS7JH3rETq2QmCpd5ndXI7Cxba
SEl3DbpSp1QEKEUaYNLfJS+PCHfQdfle8sEve7MGBqSQVrsWDxi/RIXIxj/Jj2qqLjz3UsvZdtqT
NnSfMhnexV1hRVZRKx3WGClD6riGsjLhXRvqyjQzT87wv51yVGY5C9uMu8LkWqDnSc8Inzg6TTFx
wls9I3E5IzVCN3wy+OnAduziZXxnUx0pOTGcDEz7Vo2zYYsF+uYrJm2xBh/Ge2ZpcWwYn1kLUeZV
8Qk9bR2pAgg0bZ2tZmCffnfgTpVku6opS0bTkACpq8Tg7rwzmZbMcOTHLA5lzagn2HfJFAQvSR5m
o+RAfl5Ma2oBtlVETO4GQzaIlAgULsSS53N9tRuHCqjyOX5NqMlNMlelkF3/9s8UX/jodJKFL7Yh
seaCI6Kvg8vcS9iqISKWWmNFCZdc8hrkAPDTmppL11AjjcmmKypAmRj+eVZ9ptqQNpFxUXHHujJs
pUkTSQ0RqUk+sFpgR7UzOeqkxjAOkwyedsa07NqnYY5+dbTRtARvjPNyzT+8M/brDvYlsGJ9+Sk+
h/YHLFi2XkD2lNHN+DiS/eHxYq7o4U5vAEs/spGrEtA81hk84fzriUp8hUPAQiBkseEZHQoy+pfe
yniwEH7ZEVG3fd9XugLdPxI+1y/2pJOhbhspXss0NStydqhNdkItNcobW1YHUzGVbmyIqNCrBiMQ
zxWULMKWvA0zwyGdDHWz5l36gVI0PxmNmF506nnu36FosdhDp9m4dz10R582iu1brH6FCzqt7wH+
uQP41ofefmd4VHOfDglhU/KOAk9++Q2E4GovY1ORn7AzNWdvBfqWlJdOOdicIxNCh+UjaRU/MP7p
msvXBveoYnkk3fD4GXnTuCrooK33Fa6baMkj4Lz7XFwDIiVBjbwd2kKDhdWv8UtlNBTLNfc+8AO2
8nn63LbftB3yykekr5nyMvtleEOrn7SHhwb55p3pYHdmRfCKb59gYmlGVat/6EPwXxHdzlg4Dgvy
Bil8/OUJ3VMC3nKjCtOoItZBCGzb/8U3+9KR/1TUy0vCmRAehJnIB0KAtumDIHyB6+VogBWwzUZu
7jCef1BuMRn7CjpvwkxDFvXgspGt3974OcZCCKpgie0ZGXhmkPkR0RldIB7PPlqrj4hsfuDnyQLO
HeH9CVeEWPAHJNQJ8KIPZnBNyxRBG3q/oosy4HtpdUTa8XLbGTZqfekpMKWV6LSoVEnUiuGCJ4MQ
uHnRMEMC76/N3VFaw1+OwTZ5VMc47NRZ2DXT1+ay7nxCNl52rMCAm7Mx3B9vBLfjf0UKkzbGg4nT
HioVWsN+9hoiTgiSIAfVpF6j2Zw0tyr9aFtMBmdgcxlh0Ph7uOJQ4spaQkoHAeVBE2/RxA7DBDx6
YFl2A6gY5yu7ARSsc179Kw9a3aQ5xdHSv6JIugYbX9wLE+A8eUk1GnOSYfDbRbCvTDgu/6hy6cfQ
UsNBPRu3fBBRGnx+WQ+PKuCg95onwouC3UvDWgxKZFNlXZXlwCG4uHX667Cu0NCzug0O0ZRkygMn
qsCUjgvRPOa9BDN7+bN9GiBUSLjYpBo68ibEXeC28MIPLL5az8thnHCJdl4IXq35jnsF9VGxphPA
KTmrVwe/Gwpc12TwfwgennIvjKQXtFjsIOFl1/7HOOCIwuvtVccgYXJ/Yk/DlHX+wROLR/Qkm+/2
C5quYzyqS7jZ1Vcieke6q4Q6hz0sifOMZ76fONP8V9zlw5LMAKkEebCzd/ekrAW024tOH00H7ZKm
c0f4eSxev/xNWJ6Bp9X4HqPoot+FWyARDdtRWIZNUR6fLVxgrsjkcizOsZMWK/OgIdHiFPKMs+l/
/p/4nFmmnaKGJc69XCJJLWiCfpZxz7kK3DaSmBf/UbRhEXoRWWg4iremLHUPkP7v7yWDYJ5HIkFo
Mcgf+21SwWMT3KpJMagL7fcdEgYzAEZesuefN1LVC4mbVHQVIOqGg0FvENg1HV+WirWe32/h9dos
icJTAf0ribB+TsHEjW2QICGyyvKvwGIjYTFaIzrcpdmIEPyo7jM+KetcHzYh2UYSrYnlhc2NHXck
aDi6d3EddVp0cAP2bhITMTXrhbrG1dBZ77fUbeUW0MZDPYr29UnqDdu7s5qs2Bzd7EdrxrjzdRCO
wwFjy38CJl+h8wC2zGd2MuYe3jPWad/wsJtNUEd+unDwzPjxmUDOQY6rKUhfbiyMBPV569pRSrMN
Qb97Z7WQRPz/rdlSzWS/bKpKSp+O57QimnyN9Yl7pERqlv3A8jnanbZPvu4o6m2e8PC4Y7wnEcJp
nD3JxCYiYclfCnPYLyGdbkCc9JxfN9WaSxNX7P4VAXHGspExAAgOk6Zz35XvZBFtAPMeVZxgA7gi
hVIAqQW9v9/qERFp24j97J0i+9kkptIiMx2l9iCdnF6mGYdsdXvkurvlZ9gHvRcF943lrAPqRwSs
x+J/iXqZAqPQqyrjMImPJ4QES85vXYh03H+XLvhz1COOe4CUSvRuYs6FF1IK7IvOjemlsL9Zfn0d
2W/lKZioL3ZGj0nq3M4DPYluZSfk6p2puvkx7MKbl/pp9jEbsE7S6rH/xBr3IDcFKbj+SzBLEqc/
7Wr6DCvI6dL7qD31o6IgE+zH6pDYNRpfyqfAqvvzyxCNZukTPmkS/Cj+CPXTtQPRpExp/cwymr50
hwedvTFrhq/9mntVBJaqx0YXUXnEjYj6+xm8ErMNsuPrZcwQrzndunWm77R8kqoa4VDZGXIz+PUQ
R6kBsOp0aiD/N83H7/NGO9Pk+f34ESgmkkXaMQfxkmQ+8JzBBWtiEUwWSkYtwZgkdU08zEVQVv8B
19qjMEsA1/NIegYoOQqu+26xOxsq2P7RVZJdZ8/8vgDokdCOtUQxvFGhxY0XIbDhKX85B3DExF91
rTfkhda8Hv5Cnjw1MpskoGX4ArtXz8rD1m5sLdzutvbAVDX+BUq/G3tmTnep+OjtzyRfxXCGwx65
pHh+a6JiILJLVVkhL+1/FYa3QD5uRFt9YegNrOPDLo0+/VR+IX3C7KbiJ75M5Xtbw2wMz+MytbBd
+roufZJjroU6o58wfWZA3srKjpeEtpzax3LsAWTy5EXS3CD12ntauA6luv9AdX4pktZXc/MJi5IP
4EJVKaDjwWtoBou+FBZET0m4yfskR1bf8UqwbLVxZGMH9PsIp455ZfQIQG99TDuZz1lu+/TQQSq1
3qgrl50HyFa+fc85/GEdythhTvWs3nG47WvcI/lkFqPdtrF0mhUz2fiOJdi6w2nz/g7Voo5zSeS8
rnXZZT0AAjNh5iqPJPthisBJIuiWdQC3BUjlOj0BXG9WReMQmloPH3/Hwt+k7RLt5F91VBB9ecz1
zgWRkrm+FjZmM7rzqoANvJU0CZ/Qe5367bICwyxoaNmU5yNhKj2+HVZt0hidK6soEdmLdV5vYuG0
ciEVaZyNUSI+kTH99mSOVTyxFAqrSVWDEfcl8Pj9NQ/gDHHLF+CkeV5kjcMl9IB+xHEJOuWm3+ts
caxJjOSJt6P8ajKUhdIzRR9qXTeB0T3iYNLEqGZerOK0waGOWP8wQnssyRmDkGNOAJgcMoWYbAlR
+Zz4OTHKlqd3dJJprnPJ/tYaUA/SH1Q3W7k7045R/PlvmLO6Y6qyu8FDnkfJ8PpocclO342Vl9+3
HkcypbSE8fr1R9uYC5oIGJDRi92NWiL7PSPWoEuC8/ZhxfiFs0ckj8tK44/s+nbhh9WpT4CqOmhV
XYjaEfYV8B54MHPJN1axpCDWSrJVQrkaDtTr8oWHoCaybb70InUHb59aFaY+L441cpIls0/x8Sed
wpt/W4bNw2f0vSm//cQZHDQLD4821R6U8lLlJ0MPFVpNmRs38Aygno9tKDkOQxFNbtTaJ6eWYy63
R8MsE6Ebx/wVWZQDbz19wKNU1agf3pO9YQhkgjZ19Xnm5ipExPFBgHrp6C7IJsP8qAEEiw0xJmn4
iU6BkS6VJhNRae+wFVWBdaN+WkYNr/32sZ3v3A1Z+uictL0sy2UcoSgkIsXGKZT+LHKcIiUQER86
DSI7g3/M+osmRQwoKTR6TAU8r2IfokELmGXM0tILsnrRnFplTa6g27gJC8G9ML1TRrrP8hl3Yhu9
uuwyp2aRUWK7zQ8//BJ93e/xlD6LSOa/1j2mLcGBUFzgAKN2V9Z2m/YcFZbeVPN3tUWNnMBAnFAB
KQTsXbD9Cb+VO4bPjd6XbreJiumJ2AqDNCvADIIiQq/aLL1yffqoNI7Th/jsJ8Y1kVFlK94x1Ocw
nTkCctS4nq5Cin9rVid36uv/v4/A37iM84xeVVn8ZLf+8z06EuprIu7FHoHYYMMNjdyLa7dzkfPi
8EuVgywOlsFOaKLgsyODVGXrhZL0lGwaAcAPBRRE7IQkwo4TjYbSEU7QMXus2RfTruVRIgCGDupW
v4HPtlWN5b7DhP6Zx2k+5D4wh7D0Un2v87WGw3I0CrhIBle6EtwWfN43UQsFlh0t+d5t/7zn4VIY
d1lyTGv2tH+s81E5K4pS8m2YcFDMJZxVkbU7VL4dW/63sBJCRiHbUVm5QBdMYr9Ker/TLsI4P6PP
sz0vzLXa95AFlrphp43Fd4k9AfU6/RrVJVwXR+IgAdrn0PIbaf614DoJ3gt9GN2yziuriARpYYKE
ci9lXiOxIDLSpUr8dcYMkqFjoUwMvTKOc6dKkIxRW4NrklJL0QdPTHj+qQXIdx7hDd2CZVnq7eKB
yoYX5V9CmV4ukZRXq3Nh0RQ2kH/jDevTPSDzZpoOi0eKdGrJ5kYBapzZ2HxuMNHF9d5HU3PdaG9U
8nrTOhzqHrax7mXlf9bf0KpDmj6w7cwlTfepl/giYozA0dV2juhvmi37IPvvVwU1TwRHe/MRSAVY
ZgnyxERNo2Bg+y39MuOi5FdXSwP1prqSAHUJGDxfW+8IYiVCJG6DF1p+351gJltTWUKYqrEqyOw2
ua9yuMRaFixzjXDVnV94xYZowUfFrHJytW88+nJgT+i/qkJnADDGhz1eHnZDE/XfGroXE7ap6r6w
w0CAuTW1gz7iCkXt60+2BGTQ4kvjIWX5OZ+UFF14jFPGRVg2pCzPM3qft1wXkyYUl+l7WC8iwlow
V3qBKSU3y+YauHMi2/33QCZEEHjGRJQIieHkaV8BSCSxpVekSMo0s65gvr3jbe+scGWpcdf5IKyo
p8ZacCyAU3dGVIUXMbYncq+xtTz+u2s9uNs/FeDjkbWnoGthG8G5mjrgdCohfWmxBshFzFkCKMYY
Jlc8nEQ0KHdIEwIa94YbtdIpI8PgcOzlvbkq3bmR/U8IsqZyDw3kS5dImGWEyRTpG2DbAg9j/ZYE
EqCzfSmp39iCA6OJGQYzTyQEYmDJazA+bsrRhQNav7aTU7hppZDn+GCmJeAgDDn7PwxyxdnX/NAo
FAl2YvAq7oAniHUvSxkF06h3uh4LyZJGZonVmIWWXrlaBdhdwgTqe+KS5MDZqp6+ZWKWf2Ps9lP5
KnKGpLLFGjVkj3Snum0zWWJLhvK8rRJ1qCrYgAA9OxMO2Vcsh1TGBKwz5djjlhw4kt54zGFw5Bwj
n0p/NybxTfSsl9LpyidUdhHO+Yfw58OWv0icNKwPlqnRGuhOTTd+OFRescaz0aju4/8MtfyBCwfJ
6lZpJb0TB/E19+OG+TvmNwTHUlWBEMOcYVjKqN8cisb2cwHpTQIy8ualhn/DagCriG5Ss5mbcOrD
f4o353dMOwp2gPS0Z+NJlANcu2rk3C3u+9Hic7ZkXnI2qFdU7/0tzBiHzlOSVn6thGcu/MY5KaKO
Tx2iYMrY8s4zTR1mah64Ls1K8LoJXpgFGAKij1kA4NGZXV2oHafJSyBC8OtjEEAUED7tRQU37Kli
KAEQhjAc7U+4RW2e3i0vawfHYfqYvai9FxiNfFyviQZMCrJzUuvz8/9edI7JrxdomLAcJSFqGwXf
TXosKyay7TJ6MOElFR/YqupAh2de0CZ2kgpKddDtRNzusjSGBfxQEnOjqOFSPyukfCQJH6YJDj24
wlev/3S0rJto5JvE3SxlgORvH+ZpBdU4WLZzIroFvGjUKsHFh6BhSXip914bD94KZXhm9BhmwVaI
R6ZwHDSdmstSFjgX9KyWwPSJct6v1BIhYbtD5qb37iHMZFgXJE5z6nvYh/Txr8x0K11Niv+rYS2V
fqjaSatV7K8UVsVrbB7CHEWFeLN2N5B2G2vXpE2pRZloo5Sc20AgARReXsjUfjumknHqUAmb1hN4
+aYVNJW+AbE41BW8751ZE7EpfL32BAK2A9JdtHad4xXexxgngrQ1gejDhIFBDnJ+4bjgOIwp7JR6
TQ84kIDVkgm2JP3BV5lg7zJaUE28uuBecR9sIsaxYtjj1dgAyPJnxXsRzljioQr4PmBDi8acCBZX
iWys1NvXStDTAV6pI3wUZuydvLc/oRxHLaR57MbUWDC/8pRYRJZNZzevX9uOVcn500w5rP88u4TQ
fMX6lDxVHtvzx877Pd+4Qd3/TNXvy6KHcuFOMoKl7Aw3y3G9YxHDFM1CFt82ygPn7GuXsNMMRTyl
089klR+D3UNrD4A6QW9tVp0vhx8Yet/L5uow7As9vI/F9lVL2pZ57capOWmbE00XDr4EevRizr8e
awYRcd/VePcohQPFdAdzxzLvATM9ifPFMX37vrFrs7P+XSCgUeB+FPDuApcvv9g/CtY1TFigw18C
DrIet8MznYN1/2pDHRzH6fY/uNlMeEynxoJAtN4ZoiwdfhNSszK64FqR2lF7T3c6GSpQ+BCQZNVf
KAebP+3m9w51Qa0r7XTJESwRhACxQnt8hTSpvXqBwn2KX3bxP9mjFNMKtWMNArLmULKGGCLWsXIw
Ahjh6OKF9kWvf/KrB9hVJa80pM3w5nz28S3xnB9+bX5inTpKrlmZGVTABGZQnx8xN9rAK3yNWxRl
MqMFaeyZKUuISZ+NazbMG6KUgSmcusbFEOSkyVtayJVFZDfT0c22QCAntV7YhbN6XCBHlki53EJL
YXovC6V2AO3M6WGBQaVFWg5LJ/93zdvYq5RUflLMTrR7XOUwnVqfELBQ7L2hwCSIsUzyYOlRvzhI
POVOsRhrLyLYipGPzUDYPPRfU0gODLCJz6Sfr8IstojtK21jhSaMgWjOKWZOds1Jgw3RH3W7jeQG
Jj+vUd4elJpq4OlX9wykQwg9BlXjxnDNmoWctYwW3Uy/zhK4phwgTr7Lndhb0LzHDaCETU9fNbzy
Va6kM0XoKvoR3oVzxXj6vrDRjksdG0gAvZq6+dyr/KEuWbJneLWXkre470qBwUDqEUZ7V2Q6ueR9
vG+wN3c6Mv/Q30cPnkQ309AWHa+PCvgF40MUiTvnxfKtFyMDwDj8Ac1NlzOnnT3h7WAHX1z8V7TM
L8M8fk6YExAsrz/dU+P4WKWShevTg8qxpSvWHy/FtmTUO0qKe8W7cwkYK8FSFJqZkSUR2gmvcYrx
xYU+0EOvjD+r5EbYybm9KBnBffXGhriP9LXpsNNuno3J7ipm51VsZpUqTpXZ7pRNuB1SWNYs5IrN
AZZwDUM8wEOO4IaO6LJgc7W/jieYywbyrHMoXe2kq4OatjDAzBqs4W6Q8cV1gpjYCdIdsJ36G9n+
sCWdMUjN0DMiH/tkPu9k9IuuP9+a/NIsC6BR1ZTdjA3QbRniBDJPoEJFXfvmF8uK+6QcQR9XVUG2
SimZUilAL1TKmhVYlbqfsni6RqfwFx+pzrxZPfBix++puMmKLofsb+Fwwju6wr349uRT1MEbBXIe
Axw/guRifni33vQvjD3M/k8O1VrkUzqPoPgTcrffs/AP+WH+iHHUVNtkPl769dPRHHCgbRaIDiiY
HD8t+RBytebLbNwhTzrZp58tkTY2GgZiXaroqxpPUW3tA02i6XoA6meTQ/OsekXuotw2cXMepaSd
WZaqkHHWaeHVq9GABShmwoBJIT1taHmouWHz6TkHu8LWwQ8gMguGjjCmNKvDl/tPrqy+I4rf0y3z
bw/1Z31NLoSxx3s6gx23jKmVzXSe2fQZ+P3qFpLtZ+P0f1Ko0v1SZ2+DViqw95FbSn6fNoDh3cn6
uO/6QKkrZYAo5N0S4kw3z/mHKD7A56VBF0jwTUSwMZNX8yYJ6tLskisTy50LzQMcBOVTKhuNrnbI
EIfw1c6gfwe4E984UbqlscNWkz0CxdjXwdgBkzpmaqKGwpv6TZNYWL1ynvK4gWmmkZHggdBAl1Pe
hJeoxnr9k1MJqF5o4UaIYBtq5KXaOdB6uUPymiLEjdeDKS97YagfDrPlPCXkeun4U+aWfjDCmLeQ
SquyQqScW5gKFWBnEUwCQjSHAHc24q2TLVLXbqmvHb4B+sr6JuhtNdkefLelHr74pYYu5+h30PPA
zUm/4XxX2xlut+HyBPxhUMwUSLkBfm79M+BQ8wz/7mHfs+ooFEu/1YSE0nsf+cq5DBBEb/5eDtRV
KEdytxHN5ULXKPabXHffhWtF08hxqTbOiyA0LMkBPwzxaIcUEzPuXkxR0w2aAeTWSSpTF6FbLdkp
UABH3fce3haLHuK7QiqN72JvhXet1iX6Q75CSI/U2bpnO55HAVgfMwDthms94fgUHkTewPSrkNuA
UxtRaBjg2Sv/sg1NXuOyqvFIuJtnhb74Wckh0mzshlelPalG3mVetGjY9/rZ8921eIlloIyEWS7S
w6fnIqwSw06L4zQsamKzkjXVgRiUzZjexoAwvbPTm5u4JMQs34g0dROglP3Rt7onTFKJjK122pFK
C783uyDsJuR+eyODNYNdD7g31tlf3W4Xs6hQw6tH4HJavAKTfcp35Q5ODA26tAkFyEyw69cGCYD+
qumhFhKaxIschEW1EUDifZ5cxvBrKHk8Llm/srT9HEEpfLnve+UeBlceRwDUqP2c5fOwAIwjSL+g
8G4MU0hdx6CxhprtjtWJFvc0tRjUsmrdTHJLUbGWyhgLbaIGfADPwjWvHHMgSXqPDY0lKLcIChpQ
w7BcXxACVZ6BBh8xEgfgtLYwbGnDaHDaV8gjlg2VG4V3UNX1Or9vwHXbAQUZ5C2x70nmlvtW+TN0
WnL5ytTBTnc+HFbtxkPeTJ+TmQ0gp+EAfq8HbdMHxVpBJdZN6HbgeHfJYA8TZKMYrONsw2hwV4/y
nhunnO2ZjL4H9R6f9PT2iv3yzAyGtgDF/Qa33CHPqRw5j1z95kfFEWj0eWdkiG3+4Dw5ks10vlTv
92Q4sC4FWoN57RT/kgnwzNDSsC9beoh1An5h+NNxT4fgN7LYc4UR/J6FFKUMD+XGegFs4Qm+Btoz
UHlDS3bp9equ6UogCAmrZBB8XvMOgmwWh3j0Yywjnbmqb3IyiR/bPQ5q3rLSTF1Sor+N6UUzwHiA
q/ARvgzzghi/14qQqDfSaBQs3T1ThPsec9jyBkL8KnSpPJCKhptqi+clH/VxRfCPqHc5O18TBKPT
shATTRTwyenRJSkmjYk+mDlGBdt0YfIldVEvx4hGe/ji4Q803i3lSFSPs9gi8SNzRuMnqSQeVU5W
GXzbXYvtCoSPEVPTB1kUnUk3iXEX37KkhAfa/yDhF5nMJeuxgDCgctpmv/VoJuJx7LU7YkEsxPhf
33uChmq7WPOuNvX+ZbfGTz+zLp4miXUrSztaPz82jMY7XbSlnoUMxtbAXnX9gwtIpRuR3KUlpBJH
6FznCVUe+ww0B4SPnulO7jmXPCDKuK93MXEgQH3s+sQhXtMkBUtP+rZstSG0+SaNsULuzDf+7+ah
Hq9/AZdXxE+MSvls+dJhR4+jVq8hdKKkMAc2oQkVWnsPK0P77j291n1/pn2J3A6/CksX0yqo9i3k
Baq9xvFRJT9eQ0EBzZ9rwbizYN6cgdZxiVj2iMokK1aUpvQFuiey+yL6sKR2TkspsDL5eNiVvKoG
qMFKeluF+CfTJCA7vqcVQ7SDLcoGAVJtVf+pEqe01DByqZlhDWfitKKhurkVHklakuLA6Kews19h
I50jOL8W6HtkRykVSuJxlm7rDnw28zk/H1cbR5JuyUG5r4hE05o56G0yQDZVs0qsTdi6zZKoaP7G
OBMVJs/kTUr3ecyg21X+Qq8Dp4A7zY4zzyceEWzEBYpYhCQSWyY1hydKZQ2SeOGqvWiRvIgRpgQq
yyouSep+bXI+ULaV5x+pgvF2GXZ+lFNtRP1Q68jJ3zuk/RELj2K0zVQUwI8Y/5ahDO3ashzaBrUh
u1Sava/UUET69jyc3fRQVzWvyNG9U2fYOaijaWR+r+BAx5TzvrhyBi2Y+C0AkYtbXGzLjU+U12N+
sNW6inVY2ehfD3K8zx+gXGhs0wAnt2o/yEZbKzBVUY8dYDJz++siHXnnFLwlOzpkWPLqVoc+++SC
k6mfrlI/HkTo+QZa7c+YzuaO+NiH3hg7i01u11HRCsqEqnRElFYSduNtmMp4zR81Yq69QXErG0cK
YB8xDc8r2joL9FNGWQSq4Yj0RWjzBjz2uXpoTOJZkJjtLDQVzCBIQg0Wsp+Atta+wH46TOGZp5bC
uT7+MEUXNFuRJaFbsybq4y+o1LSg8ud9b2Lkusr+HaE2Lp7M8MZpAZuzUBi3EH+/tkTX1vWDCRdD
u9H9IKTnnMBt8X14JDmPOTb6CTXq8bSWQ42F0sg+K0ukf1MQ+ImlycEcHGqFUYeM8t4py6BFhzUi
4NU/vjc4FFM9epfx4cR5uIrCIHJAxZ3DQqD8mvlerC2VIgZASodsYI9rzXUc79d5jLLgbBIu/usH
mzED1FhqLD3L0lm/wngx1budc2j0z6+JSWiAw1/UvRJZthFN0jgsxj3prDvwykdXxCgOV4ftveWq
on7Ij1YRRfeL6iY8OjcAgQGg6SIqRM5aP7SgdO0jbaGJHB8KY8iWXAl3w+GcjxH2HzH6Mh5bykEo
lkitRNHUx17cvS9nEtgj1ZNGsGJUnhFVLl4+a81PJClCnbNqDpuNwHzn/zLxMbYIZwYv4mJNAvGb
9HZrEKuw3NjB5O3dGMBlr6qdExIpJq4JWMEnrQh4R8SbX5w4EFAME8KjkCa6CdyjJ4vH40vlwHbH
qJsq/ssR4fIDSQs9MfGXY12VbXjOj62EbNYu6J1U+OVoEiCuOG97iNKw6IBia3nt8zh1br3j11Q7
1emceMZ+ACfWCbaujEWVXJW98iBOPU12atgjaHKKzNtS7UiPfPsMWa3UZy5xfH3PYJi5bcuVHu6Z
MbraRTx4BbEHwz9HZzIhu+l/onjq5LuEmb7MYCCyYCnV8rdmOLgOoQNnpND1U+Z1Yob+R6WbCI/u
0GAi8r+uf/jrwpRFdg8Fox/534LRydI4O2jWDdK/+E/nCuLtK3FgnOapSaQXDRa3D+xDK0Pp/IzG
lsH05lK+fmOh3PFYO4dvWehXcbNfDe2b3imnNV86SOn4gqsPfWl7wu0ZdW4d/5zEFZd48DpwZ/di
E5pzP8Km0ZU9BwEjf0n8ajwaDGRCvOT6ZGwcS04x0av/TWJq1SpQh5K9qzMHXAO+Al2tXPbnEAF/
pVP3KdybRBkFTfr+o1tVwLaQcZrfATBvsVSgkKR0BLVUMZf9Mir4683xwQ7ZscBqpjbpzcsGxpKl
lidB9pyQMGV1X3Yd3p3ZG+HdmeTTC8IYmrDe+yFDKV633FKvqXJY9R54RfHn2uGqkOcONvZNmJy9
dKnu73S10A8qz3OJ+8OkDHZ2AcEDax9MMqQ4pwD+lhMJ+8byiszRC7ZWx2rNIWtN9Hid6j0Q0xMV
vZrPxpnzI70PSyr3NmlFLYgt5g7w65PuMBYqpRXYD9TSgweAtJeMjbfPOgc1aK6TZQji+9P9piHL
UQ1VBmoQGeIt8PEXPp7AvIXl2JY5092cw2OanB0vpfKDQ5a3Ew6/1JqudPWEQ+w8hoz6VFSyLNNt
lzCNZwMx9vkBLmJRKaTkkWsrNjCL59yBexKZ3lKW+mTWmQRTXtM7+B8yJXjrzo8/O/6VRNcun7OS
HjAZwTp4Hzy9QYFb2NIUGO49x9lqDPsvuOAM/QBJFvKq3TNBfrbjZ8FPw/e1GZkqjjtPPCKWxh/J
BZFDrbREXUxBl2QP/K04rpduF2ejG9ffElcAQh6uHYSeKuwtYdLJFf1nG90ILrFZj2hJwbUbdy/q
iDlZix8aOyvZ+wk4Al7PwRDwt3FqZ0tEV8tPyZ9h6wXnMe/sAfhEt0+uBMtQJdFwHQXi3PhKYfm1
ljirOFoDy9hsV3Ysq7TXzTeaLGd73TBPQVwhM7oAs7u7XU1P5pHB9x4xYZ16V1xBUJG4bfNW3v1p
6KRH3ItMKDWghIOAy9hH+S8pR5lDp6MgrGZZOqJTVJfBtrtiS6A474AN9kVXQ20qgpMJaxSChNzz
t6JyQ6IOaFEsKdKF0WWveDrcYlewiHqq+AXYGfN+2izf0Tg4gkUK38EFttRw1jtrk1SDq/y4nt2t
IHJlsRn+71zTzk2/57/GPMifoJNPwlf1JruWTIqsVhPLF9BAEnxnlUOtDzf/6rc6ylJ8iUeY0gMW
h8VRJq/I1pyZat2akPnhBII71omioFUo8OdR7RU2jAuS4WCSxgZz/9U4/l5xTEPrhmttMZBzF2Kn
MU9UKMP/BenYTRZV+pE8Fmeq7uTDBOScIoHSgi5PmcMweStD3mJqZWqPeXqKyYbkRBtCBjOX3Wcp
Eu/y08Br2ePaKsyadj1Lhy3rL35e58FAZ8JRlCaUI1UwI2N8Ebub6b7RMAcevD9V1wg9HtlWTcEr
kyIdW8aRjGHa6cSvW+EgC+dvA1sYLJDX4KFWOJow59G5G4pTKoGsOBRHoqmWKaLv7AYjTR1dd+6c
gz/Lz6x18JL/1N4QXtyEZkO//G1rw3RmJjvrs2GsrUJWrXBHCCsxoZK8yeYuuVUh/O+DHNazTZP0
kLacnfpOGJPplBFQSbANuYd/o8loJaZIvKLDqaWNKahTz6v7ORJGhLz7mGOLzXNgJzKAV8Rnatex
/jbV/hG8iSkkt6oiTvI+dagGiVMfnx11ZEPh4AMLGlr5fq2Taes3xttYXFNNw3rM68A7PD2q0AcK
RSr4w7OIRxNfr6gOzhxj76HJrkh4v7Ub9QGq2WWzg5IlS4OoFGFUHDUZeXKuWkrVw5ZUOJTqF9Xo
SUpkR/tN+ys37DoUMs1lAogKWkROaGXmfgYnvEQEzgVATpJAPTVwqG8hsWFP4av0/9VyUAoey95k
GEsJpwAFx34eveUnherm+w5PL5M1rCF9SZtOLEgTvoM0z1RA68oKc0/9+aEjgaEVNkme8lX6nAWZ
9u86NMkDj+zm74HtHMUPsq33Y/xwKHpPDsxmhqzAGyRcl5xVdBLy41aD1EVYUtB7949yGYOHEJaG
GgePu1Wp1K8TRmtFKCjJRK+gDL0N57ibj9CdHQMuC51HZleCjCkzNLvUEYnisB6t8YL9Sk/3+1FG
Yez6bPREl9PGlFGaxV+egk9de+DP1EexLwC8gBNyB2KvQvNBoFZ2+JEXSfJENwc+MP+Uz+Xl4wnJ
eTUIuqp9xOwvbdpTKxE9XCxS95mT5/UAH/35/UJzX/gimQPULJ7oCJc8lYditIKH5xn3ylnzEDq7
QvyXhRcCM7vV8qdqsHtzQPut4n7G7AAyIDOsd5CEO0Zqnu+zZk4O1qL7/P2tzMnB1LgIQNqbsURb
Vdd7ZOiE7D8/EGd29LRTC91Wk8NAz5U9/g4/pGKJLtmSvW9LUURdm5oD88rBugd7zRvhhFisbGcB
fZDjwBO2kYAbWy6r4ue15wbN3Gw1JnD8hlPYkK4GJ747Dym5Kapv+zfK6qQkGoJsLTs3G6nnqwYV
liymxQjLOrHOfpW9Wuti9n0Hay5FdiflCXZURC/lxeyFW4GUQCxC6wpk5fIKPIedzLBwmuA/icMT
wzGMjRlWPcl8l2Xik0wNSIp0iAlwCEhwFX9nXP8o9JUR47ZKuV6KfXDWeXL5yoLaX4Eom+rOmsW9
5u6u8UVmEmzaCrSR7zIqhRyPQipnVfixH9FtQEzGkhhT9CZeMOmFMjmuoE6gSTqPQCb+BDEj1133
6I2YeNqGW6UbkZYlU1ePBXi/RPXnd4eJV8TKFxrJ67N7r+7ndmS0wIGMGvCgSSNJeDO0hZLWWaZu
GkhPAUDT8rUPT8tR6fDMRksNbBVjtj43RoN4f+uyexnAMfp8oqYLdtHH+p1zTgH9UNDK50d645VP
cYSDnoe3QjDYeoXBWU9yU35Ci6Nh31kkrLOhccdub+48sxvaQ1WVYeztdpTjY4jckmWqkEpheUO0
2eFXANVoLaWRwVtKZRN3qEf+qL6Vb7t2Eyjrz93kP5bDggpKvjOXKfvbbMQBN5JP/sgLYbbbQHcT
oLf8sJpme3S7g+WuEELl/Aycl10oV4c2VeOpQMGTHaMyhz8LolmEYnaJsk9+Gk+LwRc6ATCCki6O
ZtQIZUSp0nPzM/yBnJgqEvvqW0rZmc3uCoMBTpZu8xE4w+URdgbs594pv8ahtpIWXmu9IYCF4tTs
sU9EByPrg+tHAADjU1Coa1WdK6iaFj9DTciMD9fc1EsKNPQSVB377sxR6OTRatfXzdcSxXwIelk1
BkRC0GA7j32ERVp6W/Ur1CFWCgNh5wCezzkT4EZ4u+xtuR2O6qzcTM9Fd1xBcBFzOllh25ub+YQ6
7ORoqb0piVIpi5V4Exk4iOZbYvyv2+iw0Bff3es3RmkskIJGuBilemxhooajp27jOqrzY1GBDIHt
ahbKUWOLBS2gHfR8r6AhkFoSonyKpjE/ByjKRbwUQHDksSKWhQ5ExU1HT55u7bA+/MfFHPQCluRW
Qjt/jRc2CLg7pSgst06/1y6QtmQ5Dg++7k06tb4ew2Y53d3VtSZ9oJITVFsl7EkdhNwrhBl4nkr2
Bk9uLrW22Vwv44Ok+JjWCKP7e6PCbTTCK+KPSiPF9hNk5YK4NKYu5fv68vLH4MsFz63nk4CBB4FN
C7w7Q9GsRZsCiFIo3kvTCLxfju9WRXa3eV1psfDYupFrEOVJwUDFpOGp7MUl3+dEBReudtCtXJ5s
e6LOLElfGByQ5V6q29tJFy6El7LWPUCSo4rSE4tWlDnCF+5hoCQbLZUmxwIMnt8QmWlUcEj2yFH/
Wvi7qa4hBAmKzdm2VXwKiubzhmbJKVeGbfkpR63GOxO7ONmBZWR6UR9oMMXYfx5slOZiEcsdns7f
zdrmJFuEP9ZLSwfOP5QNlYNjiQfIii1LfWXI3at3T3Ic7j1Dqz3m6q4wWYkydeUHVmV8BxaYLu98
2oDrcLia0N+N7akNaCcid0ZnYgdQsLDWtAYJTlqO6cJBH8ervwqr/Y9snkRif2euBRzlYtmOwXRf
UQlchie/VXa76VBa+ENg29g8utsSaOi3rkaPuz0bGnrOmGCu/o+2EVkczmLsuL1BBXH7nmKkKgjm
fMqg6uH41vS5JwFWHpGE0pK1LyWbeJIvlsAsX1VfYgeTGRbl0ONLZwd9STBlu3xeA5OiorI20oZ3
6kyYN1W8hDgi0zC3IiX/vhGcF7B2Gv6/UqylY/Z87N+uXwYwsZsteeXqquFeYQV5aZwZxBwDcAk4
61hWsbEv+xCi9cjbLW3aW9fDCeIjViQrHj0ecLKMB/VhfP5OIbvufEvg3NWH/u8m/oy5tWX2naa0
7IgaKAbBhvMgCCUeyyjYPvjxqOzQtaaHE5e9QGkFODikUGpT78WBoHA5NXGVD/8axDR1b7/b6f3i
m/+DM4VcPgDXg/eqJNcinBxbZVTfVZGxRcTf9P3wmxomCJ00lr3fsdiAbPJ7VffnTvR3QItOxd1/
N+z3bwsVHt+f4YeiXSFNzl5t/L/YUE0XNPIBbt+bcIxsiRHPI0Q8aH9NHaD0JjphjhZJGN7FM8zr
e37dwK+d6Tn4oc6IpkNHvRkDBpJpNmBqcKr+d8310IIkmWdErGSOHFHa0wejz0OgL68kHZgD8/s9
Qa9+BoVipNkYvu5qnLfNjUEP6eGCxTg46y7UUtlsaMm+WgqlMVHXNKCEwudLtzmRtopu7a3L+2QO
WLTU6G+3E/I9HL276koxwob4JYqzwJptIxljluITOku1EIhX24ijm9GDioafBVMxaOX3UQO3WAiW
rtnR5CSRzIJkMO2PbFkcRUT7JLhqSmnk44QiBQng04zYNgf6jrv4z0A6n5BEEeO+4fEcOabWM86a
wglZ/jvps2///eAd6Yx71iV5PLwE0icOLhHu4MvXfqcX47vXcqJZvj1T0bZd//LVco+HKkS4stp2
W48rqVyiMxzfZYYkPbctKuXHweUP/Fy/DYMlio1nViL1mX0T8NxrTWZROAWZs/4Os+l9G5v0TSPs
vuCuNTsCG3Kz5VnQR+7uoqQo/e3myStN2RlWP4jqajUz/vA6x0j2Xy/MZTxBUSTNgUBYFsazRifM
3Sx0+jnAOfU2JDY/hg0D6gXPGx/IBTLvDbCmKlXP6gpWH9ui7OuL0Ev4UcJ4/UHA7USF57eCMEOt
d6i9xWsFHebvJuPZyHFDXAxar+NXs5aJ9kYisFQaFnmSxwv+feGhRC+DXp8qBdgfUZzu19Ve9Yag
SyrSSllY6dRLxgHUlrdleo2+rs6GagMVNImigBqDgF/wY1obC/7Ohsp/V26VWbvKXHFHJQglqMcM
tNYi6/Y4dMbRQB0fM2dW72v28ECYxkisdYOl9CjAVWGxVaBjew8IjFaPW6WT0BNQ3hzLYFtDps44
ifCBQB49eBvL03WAbBFfZMMi4WrN5cbWel0OsMXKz6vFQ+ePWtF3o3PF3ty054PXdVY+4tfk+tfl
uyUUb+auteCi8kg269HwDPFPqN16dyK227dE4nRDdAnC44VO5cOtlaFmMsQW9AdnU3KOmcS04+Ep
Sz4RRezwjv9pcc2+Rk25ixFxP4bssKDfk1E5sD+ZnzjYc5huiGKH4BhushPe7/+yjc4fxeXhE6E6
GKOCX31ye3VKG+bHBQ2j8rhy1Y9AQ96CI1n7H0gOXP8zx1QWUyOu+akXx3oYPQtjPHmjRATAQV++
M9KOQgQiWdTySoosJViFdEb5jFHm0cTswtEy9ZiGxWvjfRKpDozrLf7W8EzXBBTpm7PoiBX2cmo+
ZL+e95pjTUSHY9ePq4mFMpX0Ylrji6XzVzr5eFN++m0s3XW5C+U7lgoeP63OZ81kMxramkpyjUTA
F+e1oWBYX/i5XK2wbp+5mAh5fj9EgVd2/+S8TwwbaxZ7/J+07DhFbeCW6xZy7Yrim00OAQA8EdFt
6lTfGasjJ6aVauqgZuCGyD0dpPjyjtm5EItjYFazDSYIVc7W5deJPMkz+LBinG+/58kIDad/Q49V
Z8ckRdVZbyqeyqcUa3TqrTIN7hrg8WT6CmdCtxwMt8HJVxjvy8oEHeIXWC43tqT/Mqdrw3ZP+d+G
3jPzIpoQIyRaD+hhJfai1Oqaq9zyPSC/6pfGBJRI5OwnDZ9ctsgHeZ6V+/WSRiTwlSIB2OyCAsS9
rkPZGEbdwWN8EX03cS4Ov5RQ/bS21UP948cRyNsSBQCZQ0fZ+QS8SV5hzRUjUApQUb8RYbeubzNY
jwZL0m8/rQp9u0inFnqpqSHeK7O9erbVxFC3ZhNzxjKbYzzdmVC+FosTMdDzLXtOreNcwbDecmDR
/5NC9aflfMyGO8ZUippWlK8mnWO8gQ9EKbqYGNjWt00vDYDv9yZfwR4TqaQPPkQY3inahsJ394Om
ndnrv0SP8NEaAqXupGx8OPATqimOr4jxNCSBNrLmb3KsBUUDBDvRdYfc0/kEyqdTuDyHA1ds7Yjv
T6OTivpY4NqnVB8KbNCLYNL5N7j3JZX5qycFKMsEo8XGPWeWOquPCImsrLWZdaTJ/I2+JtGZqFLN
YcS8XHavU8sBq6XOwfDC/zaU1OwAXdbZvk3BvXJAxvMr/HKLWvJv/wmEbuBZAkb3wU7rHEznLODo
GHW8KgFpCbofp4EJ6ebzlm8h8ozWmnZ/JjjVCZ6n6+0icelsCyl5srQPDqWBkuaNSlr/ubf1x8+g
XZnbdCw4U2ObBRZB/gFKWTPMo+tLPIyDXgoiW8UfYRXb95n3sVxjjT3L/IYCl8Woc+OD9Sh1Ibes
IvkWhmxgGyxuZ8jHcf8B43q+0gqyliAZx7oj55epElEfe+sEyC3SPaP7TjkEHkbOp05R9lKlWKNX
VQuFzYVgeKI1hmUe0XzGWfY9+WmYdJPms3FdaBIMG9aJD0TjA5pZydX7dZl427aXUF+XtkbBUrRJ
g9o6WHYlsN4oOtwNRgVlja+Qwo1GahilHpZOZOLYvx2n3NJcVaA8UYsjVNS7eRXfX+P3y8bHSgLN
NFNXwN4SMmA8FDfaKajxcrIh4r+IxzC/Pjk2xmWhXptkgITGhtF0F9SrAD90g/7ux/DSzh9cn4ov
qJevWtQTk1ugQLvOZHQ0N9l0fSMe08LyGnLhWQFYtj0Cw8BclmcJTodnXHp0D12b6r3MEMCvr/el
nHe9Ibk1x1HwOk3m0+3nI0Q1vRe7R6yp0weCr7utCfEe7jTiZa31Sy2OphOfahSDeVdPoEl2t9tW
SdJ+byvwBHEWdGgMDQnVIOHEvKNyd8L0lOmtljs9OK2RJcXluyoTaYLiU7ldUtPryXQCE1HtIeuD
cj2e4TdvOSRflQR2nqRayiD3Vx1sgPEubQzEFK2lDt1VlaUfWrNgUJp3ULpMd3V6kwEuSGu4k6fi
6viHxgQFMY7eOwLeWyOc6j+4doqk6bOXh0NHX5ZKtu6bnAWQIjKPs7sWm3YfcAFfT6eG+hIagMis
gB5oz9CYfWo8HnNxz9qV9AX0FZltZdBEsBcSvpbn/ggoPHLfw/5nLv7snyTXXFVKlDJmIve3LVkN
1h74RaIaXxiDWYEgsnU9K5Nf51y7h4CDaRB9ZsDoYVGNp68YYoF8gUGrHY+1Id9FsDAS2gFBwZ5e
4nMb3dRSt+/OkiJvknD9QpsFCFivnu8Y/vbCT+Ydh1MkUQooutjvhmraK0fFgmv69Q8deg7ed6q8
Ui62eKVJidAlJDSqOCiT4dig61LN8gCb7Yf0WM/HapIUjQPAn2xfyEV98PXqnGI6YeT/ufmpeyV9
5l0LTXQZHwLummXWaHP4L4b0tTxAhHdDS/0c9BgBcnQxzCGgKwfH4UW49FjjmHBne73rTQ4opgTE
BlXJOCpMDZLYqc7R/UCvJckuZHdCEmR2AgZ5NNtdghP8qqumd5Atw/Mz2EQnQaqvk/42ldVFuQv0
OIr5TeJdnYU9j0AQniU1HJs7hofk/M4g1M2FZjWZUvkvMwXopOTtkG4KsykJ2la1ZlpE862UOZSr
cpW4Jpd1AU0Eoazl1lKuQZIYxUQB3laqiMlLt0x0ZKiq84hGjVu3X3VaZzvg8NoZFXsBcp8ou16j
bhfR7zMdrKkmrMGnnz94r9JtWJ7Sy9hDRtVLtcYOL+X3yQDyMAUM5ma7zXcfnUG2gaaOnsTMwSwy
P60BH0vOOC3R5J2oj+Q8BQ/FF26FZZ6NHioZBkOyqT5UtbBJBzueVYViEeIZr//XRB3h5B6riDvf
O+TR4TYx0MrSjyIKMLsNKGvrGJQGM5uIi5d6lOQ5N8SFGuX/Gz5sSk1No4lLOMpgDy2AJFscKtds
MG7pNBoTigsbaNLJuOuM9WxWUktSo/6PNwrGXDOka9jm2BwVxzc1Y1JAOtd7cHufpbNkMq6mAPtD
G1Ni4QoZA9U+/4/ZoxeTU9ml1ytgeByRlDFyBXTdSwwrQx701rKYQXPzLniA/mvCN6eM9qYxNI3F
txhATsMEgDgGl/gEfvMsXjdtVPZ6UEYu/+EpveoXdt72MyVIjfROyISafK67mJZdPKSTrnx3gESi
wK7Ra6VhVJwJawSDdSXsgRaDYhz1q+IdJy7MRqbMj0a8sWaB62w4KuwqscHSv6FzGXsoXGu+OaeJ
VZpCFA4NI6W0fYg7nM1BjJqkdP06fhBoxC52WpgP5oH0UDECEOrKqgyXdqXwhZzk7/IadnWkwM6n
1CoF8IwGa6kOH2WFBvji3xGepHr6IKPv7mwVeKtIEF9XdHuhpJws9S6JeUoBVD6NZQ03UX6A750c
GtHUbsjyj9Un/t9XCjQdXEcxjgyyrV2VSzkujddjSZLPqPhUPz1xirTwkd9EsrRVnwPHB1X0JmN8
p4QcsmOtpd5Hn/nblS2YPUmiZbNVw1toMzQ2doD5oZubo3G4C05qW7aiOvAwXOkVmVpEDA/OWt9r
yKBZ5J5uIjEnFCHNNNe5J+wo/dtJuBO+7qCfvZQN1u/7uifModc2dMs0Ff2Ge064IVvd6RWWOWsD
POTX3tOLbKRi1sb0zNq2zJswAywZE9f8UK4QPBF6NkjFF2tFoaHu5pbks9h1rFsVIDYBVL8hNXN+
ZvUEoGb7krv7VQ6LwjGyh6+Fr5qOSmeGpU2nUhJcRdW0nqbznybaCJVFVU7buENQdHR+mMJMvxJF
xmYIwWu+y/O06QrQ7PI6P8+sOhL9dtQbBNTopEcAxKje9gFwDoMW6OPHDjnQe9C/BfAZTgqsO31J
DToKmDnoFWoO2JmGcIOnLGcmD/R96vJAZUeN+6WeQe604FbnoDbr7Vn7ORa5D/RuOIkAgjE2flJY
dsPIcNnMjkZUC2rr5YvafMWnZU3RWJ2ItLmhjyW0GGpJKy7xVd3zseBCklac/aimycZc2tnIajFy
sguzAx5UkwKM76+Nm4RKb1vZasxuEIl3dnFVYHC7Fb1f9I4S9AID1mzdh/ADFn+XIspEHzMEWdyB
Yj9519hgwnF2pXUoC4zovN2PCDMqFn/+LuafL3L97dpea6n6X2fjPh/aSdeddxQXGiTtE2l6Z4W4
9Qka81k6f4o9D+6fw8Br4j9f5YV7ncxsggsBIguGcqweldLoLQpa+ivjM84NO4qCBxO9a5rw2uKP
pNz0R+7Dq5ABmCAMA/Ntsgy1IAskY+qtWrP2oN5k7qNWZc5ZQ4k3mWHAf4qY6/SXBwRiFYVHKUe1
F1oQ81xqGH8bPY3cnvEoWWt/v1U4bst85fs97d+/VONQXTnU7+CH07+Z1nEDX4rKiaE4QfUMFirN
dL/qHt2oUdgio4cXDeDVeGakA0Bm25RY3WnUejt0uJgC4p1GL3MpJaR0ourHd8cCbmOf83jltNz1
GYESQqflw4r5EO0ua6Dj41Xm/DcyKscmbz3K1OP6JtBVXKusc3XkX/ePtugKERQTIdXJ/rCpc3ai
wRjT9FeGDUkFzlvDoaMRm2Fhi/to9BTB5LbyDZcmeQ5TF+mgz+FzxmJ4GjoTGdMeBIjyt8e+m75n
ZlvHH3dXSOgkhR/I32DtUZ16Go3E8td3W1sKIS1LSntJ0IfgJmllVsFiYppsKxzy4W9DrcMxFPao
sHKcRFyYQZ+Wgl8xwF0W97vbiVwsezF8l+qxbOwDej+l0hs02zhOC/A3b2AWQtxd/9ZEx/fyQCkC
F/tpKem5jITcjoou5Xe4safTH5LPGIMsG4GxaxgnwW1wxZo3JBU4+MI4I8OBcz515UHl7j4+qxtI
48LI7LPE5pmWpuvJYCpdvD6KKSzwFXuMtZubJbb966bR96Hp/RnCxLPAGnLm+tLzBricDmsRILqo
+VV67Dn3UsELjXpnjMZQb9YsmyFOiopdGNPuieWbfcWOsQQ1kA8XnXqTolziFaUe6XodpmCeKebq
RAuHwBruNMkeKxaGZzrKdJuEeWfzeeQr/1M4cf1L+dGfUkTRpvs7gGjgJl2ah5eiuTHZNrLo7ZKM
WLGvD6NF+RXHL6uORbE1Cru5KLdKF6jIS3Ue4Rc/OI+AX/ui61hW7qWct0AR/RLixq/MMGPR7pR3
xw1UsTVsM42LdcqRKQgMX/buX3DCY644RfbEcZaOv823UpO+aiu2H7fFhPi3IyN3rGp5SJ+uBpTG
0YFK1KXXnNFNGltJ4exLnEyb86GsJxBCnkhdoGLR2Dlopzp30czgMlyK84vABhw0TRDTPLtnNgtc
WXHgxI+Po1UockurydlDMOOscsW9+KxWvXlzxa4D2NVzmik2nzWAHA92mR53zUhkvYA7ABvdLvoT
+7rAL5i+EmK7JXMtREMnSTnlCh6YPQ39kfpgqPSZK/C0dlvlBKegMh+mu8ZJ9rE8JYBj2my9uGD9
tUP94BnGVozIEDsdUVsFhkecWExzm0Gfmo6JtpIZVkd9SF5TzmjlXp+ShWmW553NWX/byPAD0GX5
tNAalEk/IaQYjfK9fQQrHuEAEBmnNETNHTNOfYsMAuNYb5qTsDMNgIDPV3n64SNvTw8r1tgf2MlV
nEWDLW+VTSCNyUsh4kvySmG8zsQv3p7CPgpRvz755Fhw/8nfQfD1NuXuVsp9ZuURlGBSQhIpC3zM
zQhDJeRAUww+X5YtinEAe3swxLbD6EfaXkku7iqp/ejXXXpcmB4DC8lGy6DoSesJXSYyMqqP1uFZ
B+6rsdtUqO5MAZCLyX5LS0ul3o4KtpmXjF4Zrf9phMnfkVgZ+yd8PWrFlzGbDF32eUP7mfxoT1La
h41CWQCK94nLuYin3UieD5NLVr/+LqQbQM93Ch1oa1B2De4CIEw2hWuk0A8z0z9yGEDupdK53UaR
x8bEgALBxP6V1xwzBOFU6W9SSBqdFDOAejj5TyM+TprWp/1rOJQwJlFOeMsAp4IsZlMeKqFVjl4d
sCrzI4qEZpJ2PlK+ofrjXh1qAa7uKDUdFsphQDYfvA9tV1O1fLBJoSZr0zuaSOVJF1vc1kCrw9cv
FJIq7OK+/0+O3B/iGsA3E5yJYB+mpe8JLMrZ4uAi63orWovYzxKP5vO2IebWqZtk3F9Mxd5EXf63
bMufGetqCvaS70DVVYQdLxHhV+N4qlER5VGTdlDayPvOvxg4GUHox6zxRfQWTB/G41PqVI6f19Eb
a8PDkjvnqOS2Zd5QhLXlYFKdhqVEiVGjBU3GBPHXT7me2xKvfNdgjI+AwKtXXFaUp0BLwFiySJvf
NGYk/ke64H7yNLPf5e2YfsShhECcQaENYMrMs467J7/QiAcaZVwPt2iHLxeYOT9y6vAAkSTyObIz
SOAyWa5TJnvKLsO6mF91SRPb9ShBGK5S1xxq7iOMSXeeqKKi7hpkgDXVcyQlaF+/U3LeTwSdBolV
0OIP9BA/uXqMMZ8QT38Csagq3jQRDiyk4txPC/D9A0G64eP1PBeTAO/uwESfK0BXxhtU6rC+7dPA
TisNvXKGs9ryiZXwK6IGVS31eQMy9J/jvYd7W3pAGTXG9mqDMwEtVXwIoJcfSDQfsC+d5EsdCQQH
SzQ12wp4Db2vrdtZXFXFPZBF/T1oYCXsQhtO0ivwkSo5CTdx4HQIKtfgxjUXgKNj6/BcUF6uSc9Q
Lkpkll+8ruORIR9MHTkrdG9HyYKeVs9YBiH973g1T3Tch/ssIEi4RZdhNiw38ZlSVKelQyUH/tdK
zklg+/wYSdgbcsRxfKvmzbfhwXnO5qjdewZ53720naIS8znFpjOf0pNE5v92cKCrtsTqraZd2Gpl
h+7kSavMmjqM8ZxPhH7ZJxH8/GDwdTa7RI8QghgC1GdUN9cbzlcJKIVmR19Xk17B6ukMMcm7sQIo
WFhxCDOw2hg5KVnoNhhYmAF7iyu3ZA+7naqrqRxmwCcYf4DcSLPWp8CHW6uPW+3gqEcTg3qrGj2E
tsRJdn5JuORr0lwl0KCZJLCJdGQdndk41WMWYv8aGNBT7A7suFblRHLpb9pBzI3fCCcHn/HzIO+w
U+SFhZaSfuGUGEaGzfLfGkhii63SuSY7mn8MgJ6flqPxW43KGwVnB8DqbanQ2LgnA1IgvMGKlEdA
hRGQGIsBg/8wvKaDUcRg51Oxvuy69OfpGR1PkQyO0NaKmyJiknVvdJLHe1doXQLieehrZEqCGimf
WXJvaVXO8Ubkya1cAJEWisYu9cbyFZymOyGl4pNn26zF/XsOtWn66JtCvaOVG+UVu/yFCV3tbxMQ
rieRcVtxayLwHx+ueH469LgtxodQxGiZxpu2RWQCqXc3ZlcYEStwi5ft3k6jF0vWK+saGsLIR/c6
w6povRKSzpHOyZTR60ult6Sr3NIXn5Na27LqWCMnwy+M9ywXeUkIXUs8wvuXqLMSAYwJFf7Rwioa
h3ybDJkTUY1rAxw8ZGlsn9sU/VwyOZ6Fg0ZXa5vsJj1ay/8knHQ5Q9huXcQXPo11xX0PTLcUrV5H
AFksMpDrq4p+tBcEjNZue8s2PaR5K/YjQ9qAIo01dPxXa8pZli6bO8IjEiibmYfWaQL9eDjhhyzJ
EnJgV9y5UE/TZI0tup4W02KjyMNket4kisXfWz++nhEScrjvkK0tGdh9HOp4eJYzkDHmY1ABDgUr
3i94juoYMDKfKaatqv131pPTGRhFktqqii/r6cvzeKCoO2pHKaHug+uZ/XW1UIUZw+GE8Rw3aDoe
DKTBuDTm2a5Npxmq8MydDAAMliFp1t6osrUA+n1GtJ9sfLqP4XMXjKFZ+s7tHOaJOVIl0mqUuPKX
LEr2R+WnxmBJPEUJ8DOAQmTjn7YsP67sjh+qlWsRaCcxeR4FuwDAQ8Wbv5yUyEHkPyKc9tugdJPw
ePfXoGfwNvCTr32CYk4hlwukWUBRTVlc+nGHu8RNcY3So1Pvagu6AZ+vAIZe9TEYDNYGcp+3VvLj
80y+R11jna/qOnROWG69xIJzylY2GbvsTwCLdBvWaNAbeNC7a6BG6Hev4rPmdNxJFFfsFwVr4o9b
cAifUSdpiOW9lvpS85jKXKyU8dm+bNpha21RfxaVBvE3+AYGwxIzioPSwdeg07uZC6r1/pG4llUf
nhRu4hJwmb0Q0a9k0kAun4zySjcdAIJc1hdhPaWX6EcHNXlag5gSEAYM+odhGAS8WiLoIWhCfWJL
W6r9hv3NoZikusBDLp3EzRABPXMWhTZXRVgrJ+fF4T1AJ7C0a2p/BXwGSD2omolKVCia+HvvJgiY
RRtj4hvU9NX6BWsd9+VOhjltDltvlDcL65TRXW9rM0lh6G8SIAKvVlQ6NPRtg8IDokyNlZy2XTQ6
BQByvLfCeFUOz6jmsbkaGGUt1DjMmX15lD3ePA3/ivu0gPZT1hMyVNP72m2yWnr0uifQJVacOpWi
p20uCCxE0nxQxNI9AmhBcx7JlWvwgzmTSDnBFuSj7JU9qhAUTxPhDWPE0/qHmb8/8MwN36fioWHw
PE0MYDsNY5UP+J4ZNaqV3bch2HqrpPh2NeIotW9Hz++/iWTyA0VSSRxazoFLuTcYFg0AxvduJq6f
QwSQgZnwE8tA/1jXviSs4+hOWGiDNJZdNrEuc5JC6JdCw5sqQKwWZvsW7pHiYXF+YHLFvJj1QFFQ
VxC2lFDMHKH/uli26xMzTqaY6WbOLkNeeTqVABjX3rdiJButbJuk7KNymNa6cPRbz2tOhiSstXso
nw1SxhGXcu0lRKQpJ9V1U3W5y3Jci+gg7VZ4aTV+NZOPlEgfz60E0Etz7ymPrkbLSxFRXrap73S8
AJI+Pf6qL1kNmMMSM6r6jb7PIL3pZChfYxgIxjT0Jz39suHEGUNncFT1G6x0cfrGMqy5I5Zsc55O
tDnHCx3QP1THvT8I5oOi8o/NJ4HS9eUACBdQzWi7CLNiyaS29/qoBUHCfiCjErV27CaWFLoVpCnF
rgxtrceHR8fgvFIx2w22bTC+x5hnpcoykG5ZohBGlr76Fgnpoz1D7I7d6miJXkyFNYbmQYMpyfBm
v6Jv/B/GxtyOcR0UUeum2ap3gagFaPqeAyPOqJRwKpVJ5v4SkTlHelPDKcEIS/4XmFQ5dng0RBBm
IdBN2eO7qSLbD5UGPtUn3vnTo8rTCZuDk+6FdZucjBRSh1EwJ8LuPraAXJmJVBJvkWhh1R1Fh6JP
o7AoPw//uRazKttWB9VgEyVd7XVuA7Ig51HlBM8D2+l1AqIJmFFZKaaWC+N/CLBHFjoAZT4mzg6w
Sh/YqQCXKUIrDDDdfvu65swDLf9SopkURhi72DYNeIA89Q3+bW7DCaugOfKPItgjlgbeLZH+F2ry
u3vkGclbVFCRHR1NO4F/BZInHdJPdN1VoMNlaPDjNfkftCQK91wHKwEbjc6N1wfnEQe/5pJjDuIh
M9W9WLJIgs1B7P5bKzNtipLWbIHTdC43cALr8VMGIRXkT31EwzxBiFcQWhBk5rPbF1WjbCjfR/DI
DSFnWL27hc5Qh9KEuw5e0k+IyAeo5fPTwz8HlKydVDlrG3bXeNZoCfvZK3c7d9aWRKkKnxnto6s/
6DohFnSZkrUi8vbYsd1+UsQdzTJgxZ1p/XPdkHhFRw7KxCZxRLUSPUgK/6aUkubGe/zI2VOUCETD
4eoffK0n4tN/qrpi/opZL8fWy6VUxPjWVaIN5f4Qnxdw1+d7jyAV+sysYQHkqxPX2TnaEHQg2vMG
1FGpNIPURHZDuXeep0q2R04GUOsVCoFwNo4a5sXlxoz7ckXzEKBmQxgFkLt/eiUy06DTqu9O2nUZ
eITFmGBAdCjMlgVVuXUzxGKUNDaFWW99n9P1dk/dXZLhhJWYtftdjtMqews7IL0kNfijtzb+ycid
2IxPqtvZtVt7INeJSHHMh+WTvLejH6FR0+txrURLq72wDHlUeE+fPN6Fw+YajGcHa6/UGMfvfN5A
UvpdZyU+AfC/2+DZrjO2FK6kbGtVEHl1qGvRLjPhC8ZkwUXjWU4zZfWMVR2rHTDqi1bgG2S1aKo4
YZAqHEC9VOr652L7lIt5eRaRRFT7tD62n7QLlW5lGe2qcEqmwdwTmBiYqP2XltFz7TRg+2rBaLPA
CoNcHHRVpODEXdsCc7VbgxFh2ltymULABJMp7ELjKXvg5/hFMf820PBDCeoW29WuXSoGa/qdQ75/
QELthD20aavp5ia3FwO3ra5GTLIyi1fC4e5pxQtpIwOnYn1R+86I8LKjpwhPwvnPOyuAdwS6YghD
DsMPeC5bbQ4Kfjb7N20rQveyXAv5jq9oKIiIBOQ2vZhaA2nuTETKZA19O3yW0Q2af93VNpg5lu9x
blPNJdeOObKBlmGozb5zcPvBiqZP5DMVAhKFfRud5vobpomhqD/Mkh+Se9WLfr6eGicrUw5gWeJM
+QcooQzazCRcuw++Cdhf5F3gGZEdcys2v/WxUpg/dRgYdRG/o/hYHkL6YUeWrhcQqiRfZqVN6xSD
+tEt6AahQ1I0utdJAV3zRTAYxNKMIFt6MFgKLHn/D8EG5CGeaqZH0r+iO5thplC+mDkz5Xjx9mLL
+2nspaB8G0BWvB0kF7dVAi8kL6qgv7/0VGNLghXW+SZCs82cMQpZnIlxWiAQLq3Me0TJU0xBP8q8
YTMJ7j0pIntVqg6ak/pB6MXR0PT8xJG3oIHdYlsf/eq+IpT/hDrvIePbYOeScwc9nVcCIHxVkvo4
H7FskC1Kj4Vve/OUCoQHiChfO9ROIeu+v2HIg4aGofIeuxybRrNZf+z9b/KnMovlHIoiQiqDfhbU
YeO9p0atOPMAypmHHgy8vgAtXubmwTqZ97M4f1J6lhSIOXh7ZUpvzW+E5vhZYF18aD+u+vYOSD41
oRPrFBmOmHPqhNccYMJMqDRg1SjzloF3z+Or+48KNFF2huu15shm2Nvoq1HsaGjKCekVEOfKbW3b
0+/aFtxT4FHTG7hX92aeXdBvtG6eC6yuIwMNPIPgOfSIVAn+Qw0b6AC6CCZsPdxx8pFYrIaUWtrq
NsDerNXYuMAWHZBsxjnAH9UT59uzy6vsut1k9Ym9fjyHzKG1Fxrs5PuZr90HOQk5VKlggjjbt3Ud
+tO5BFQBU9ZUD2FBk8+WhkgDIyvKbGJDPEQ2QvU7Ae3Qhnru2GFaXl8oPPZFwHFXK2zeFlaQr/YK
FXNhqAw9kU6FfPUpZUWfAY+LEgZMakJQY1fgr6ctZRyBrIurYEezjPYQgACvSmJDoxOuk/6EA2K+
9RP5+yrc9uQdr8enAZKWkGliFP3ujkLbDYYnmeBOa1LhPh8GgP4htSlKjRDNqGo+LsfQLxcpfFY7
9VfABCf+xTaxyh0OpDfY+7gpxvDY9pNIK+KRy/B0XFNTsZkc2fVq89R5Nl0ye1UhwT80S4vVFBMx
XKFYSB/VGBHGwx2rEoTna/1Izwdj8bzBp99H2tVdfHY1uh1bXEodA178PewSWttUlcjGULWpmCMj
tQTDLlrU0Ek/9YaK9tQJmDRQTFe+wd/g24NH2+aYSt7e/JNODoaKQw7aJ+36n6u6rAgBNJ9xI6J4
rO6/7jXEFFgoMcJ0DIYTjB1Z2hi+/RiWbmTsCOe7D5FFKyPlZsy99nHTOxn9pvBZI3vlriYzOh1y
u1nn7csyG80n/MI1lfOowwiG/OGONV1nOkRUWJEWAnQNg2L0JrA0gqnKTHX+/r4zxyVOJHihTth3
EnsznfMSd+YkV0uvkI3ogon/uzSrs1kXVwCJGsVAbifAzQzM+Ri95yGs9SSyI0tlORVqj+Fzq4mE
fr6sidTDH/BcOuxh7ruRhUtaQNlq1CJYA1vNcKuWrb/Gd8sAWTbbCjhTGsrA+pa5xtaL274I8TMX
DSaIiM0xMkUPgZBy68Tkqxawyzi9ZJl1o4EFaw3fQysQ3GJd+BBttiGe1Vzl333uPFaWJ84qjKZq
UlZBf4PkQNxMQOIvf9TKOlgBYPaUtD0LPBzrM+r9F+UWtBAY7Bp7xbssgN/aNsE6WkGeoKI9QfTQ
VxEKlUuEw15ZAJ4e807/LNeVMXrdp3PwBasRYlY/7EoF5t8KhkJsabJ+mtEDzIKtME0nYuMesacx
duljCBz4xULSiv2WTEl9rI/BIB7eobW20kJ1vvcEu4b7Penga6+8LrPA7JBpxHnZ7LWsSkIghoEt
faTyQEJ2mVy30cN+KhCqqIhxGQvu0FpW3ReJioay9/DU/tnkYnyMRjQPwcskkAJVUZWW6ZNY8PUz
mDpoxSxdqIGkHVg/6sLJ8smy10doUqaXcYtYVMWmejECA1Oo+8gvRCTEzIWVGmPXSfEQiIuvmSvS
6+U7Ex72OSOWu1rahRCvRejAy4hJ0B5Xno0RyZRfLy2OI6QpCSZS2wDrTjcZrlAZOikcvyD7k20q
GsyGdhmHPd0YG7YtiZlR14yX+lj89prrsQDqHaBUwwYutmr0FN7NuXNjKEt4F4k5fTJMZD8KXLPk
c/IGATsawMV/RvKSV10iVmTflWEalwa0UOE3aSBjobGJvSBIacywcDObFTyxeof0YQH0oIIpG+4J
IiEtWPNe79RiwYOTwVUzweSmL82+r8nFaVdVgU2WcUa9uNV2w1JZdTl1r/Wj17GdiJEiR7oV2Z/k
6WwEDowHGUg8UfswieVR/ia4Xb3Tkxj0QgNusS8N+Sz7QGzxXU0qmoh6hmJ5ruwSdXVhQD+1wbWQ
sqnogdzlPESu2w1sqlYtdQmm+NQvPX4Z+OsoYeO51WXWqRqUe6snqhXMwc95agD17MG5m9pHw0MB
BYZIQj3i9nRga1FwWmJU70xRbN8vqn2PLymH5K+eKXcQl25VUc14quPAZLl/4MWRFYIXRd9YYywt
f0ixFa949j4h302rQ5qooeXRlJFk/EIi/enJGbaU19DlZNGiLtLO9BfFqclil47KpIQO5ypiGYiP
SmC/VN3iod3Gh3O5Ec6Kvv/jvTmV4wL7GmGPFiMgLD2TY+lKMDpjG3Tth/qGYdErV+pLO9fGzpAR
85It2kv/+LFwiCCIg4B5cwj9dOQBwgYEeLfrMW+CAipMcPmm+xC1P2sNFIzfSYUtc1vgc/s0iWKO
y5ALu4NWD6cwBgsrv0DNmw4iJxTpFyRcaLrvpvv1BZARf0d11qkSqsPlvgtKrvGRt+lHEzxy7XCV
dedeQzdsYBzXJoZ8K7ErprkdXeW05iPDAN37b4oHFuGpYtapzVIKQZ9offmscvdL4yqv+M98CHtF
VMemKKAaHUUr+Y3ZdsByhvDh7nG2D29Ckmm2s5Kj8Wzivo5smd5Ec+B/781xRIh9g69P4iwZw2lI
DntvxaK7fG0DkTlIRvcON7UctkOSH2sTUmzsL03CXMwWvNG4Ajz4NSlJvWTCi54aGK5EaLXZO174
SgEyA+1dQYjKLb5X8k7edKUwyp4iP7iFom4BidCAveUdkVg1aEnBk70NaaMP6NIG8BwjoPK5pMLY
aX8uwj8gPMNzfkxxRWb4H5I73YbJw1LHlBe9zCDQWHNyMDoCBUvMBnxb1GjeTjeZUITy8fI/eR/h
kuxfXran9XNXPegMVKGErgHSaSIc3smbFIgHeK8KMM04x5t5/+8E/KIbc2mH8WFMnOEoEoVgH1/U
L4n2jy8kygKlJ8Jp5zalo/tC4FYc9k9aHK9agtXZXMv+Nc5Pbd0NEsdZDaGGSBh9TgRMTw5zmdIr
l2HU2z2CvoOkeBG1YA3r0kaaCd7whL40F9PGm3YDT7evOGg2Y2pEDvdbN/ZlYXDfdjM0FcIdw6lW
a9avX4mojNWVYWX2fkegwk3es9Qg73gzXapQYJeLSP6AW8Hx5Z1B7UU65DbTnA54JRpKRVgCwBth
qJegZRhJQhRx2uq3AzaKymxqdrJWIW2n8rTmqNRYTg+P21fO99/N9QyJyyQhckl5jDOkWAnWNTye
YhJf0xTiGf5yGkn9HQW4qIA0aOO4P+AL2q6HaNF9xu7lKloXR3f/2yqkkTHEAyHs8EbVBqOyOBoK
eUfX9thqPOnbQshvbmoaUq+2pyzaLKLXR+ENnsaxe2i0a2KKey82HR475wYrTRAt7B7uQiXdFrAc
asyO8u2Qo8HeXU8NVrMXL9CSx+oGksJwXm+vgPSzCUAovNwfcXogbG3TfU9dC2UMYkqoM+06LK7R
qNROSTLqB/2E1s+XhkzLVjWW1994sSSmLom/bPp+78n1aeR8rE2UXPTBry3dGEN3Vo7xW0vZURjW
BHiHcgQRb/iW2rFAhnYnO7DcQ5XCVS+aYFHpkMTMtg9aeopCAgiuqR+P7FSd8bAoWbkPGp+y+vT5
tZF2z29R42tRNYh/uuWo0mlIoQyQSJ25EKWJI4YJQSQRH6MSFdVcS8D/c8sOCO81lMo2Bhc7ijSI
p0biN3tIIcdOoMQd3Sd4IGRmPDRJbBy4md6rVGY7b6l3R+hnBdJzIUT9l6j/AEvBa5Q0v87z0zh/
EuxUW3bFxpar/xrY1RDukQgEFw4dtzhjauvRpenGrEObyNsh6LfXBcL6Bim1xTmwzNcJU/TMhkT9
Jgp2LSTW3VsRreP6Tbit7xtz72F3lSPuGt6X7eppsF34OmiV0Qi8AbDtUuPz+V/xo+3xo9yGtPQp
wo74g+SyMbuV3qw5saAkLgU7lXYwDUzAlIHWok7W/ku/7UnYHBT04XnAhqoLn8sVRbpLXsDeD6Xg
wFIGkKJkMlaakmK7pywLNbkPDZre8zuHrL0/sI5jl1p7UVmRVjTs1nzC1IHZRftAiuAWjxzi/9OP
QV4FAMD2ZHBOPEPKc1c/DvjIwCURJ0b1Y58c+EzLnCLBaTHiC+L21yIjPP/9wmY3Ijf9zZmTn2d4
1pglX/E3l/El1GumTD5z/3Wp4li2iL/FfkPYf97XnwkuO/s88B6IXA93vR3vEZvbQLcDkKfEBQCl
L3x3hbrWHobuXRo2y32jG3i3XegBpzawIiEy1S36PAOLYqnJVXIR9aBSr/G5KzUp0W8XODpUdoIW
+iEc+k9vhp8LBHcHhvVwZLry/GfUoaSwq7gFMH2WNLCqn0U2OnU6ESwlZ6bDksBxuWuyvpzA7ooY
yEM/j3R57uffkYYVNC+YEcOORJv8t4r6QN6E3vYJz+iBBC1SCTQvfPm89EMq6tPo8IGaLbcqGm4K
aNX9hySC+WEI0Ge2iI7lSBt7y7pbWj2C6iElVNLYn8/Q60oG23PAVLVqvZHczS/rY2mYGmJNovnr
gC0jiX5Xnes70RhjvvguxcpA7AJNOm+chEzJjW5FJmtUFkoIMhMi95eWxH3SJw7/jwyMe9yUH5yO
6o3V0lRmDBFjY372dgBnPDwbgXqjwyGT2/BQAnEUMEDlkz7AKi0piGK8cfMYuOdKsj8ekT/bU2Lp
6g/nxq0zTa6hjSAc8jJWxHpDglUgdA2vXqPo9Fx7T9y5eMnVT7GozXXOmYcsr29wE13c8M1HXcir
lYNTfKrO9ECcmI8F8W+B43Vp3yuk740bLW3gVeT0OMF8um1Cby93Q7UtVSuH66GBdZVHg7iygj1u
ndVp2WZEM//Z4M9DHfKox3/FJjTqX5AtkQbVDPmPK59oqzNeWp3m6IAs/DfesrDnvbmeCbEcwtzG
iJwylXi5jK4Sx2kwKieRr6uzKd6U8Vlm+q2bX8N4roF24Y2ELvlC37XqoBk27/E77Bhx740Eq0pJ
9dTja0mxwf10HDdJ93w9nR1VHYwLML71/lLdC8B2kAEQ/4KekZm2tQaMtBa9m0hcAv3GIoVMHBSG
mXbpkw805ApTBGljOC38tu2cAjwlBVjmOrAuRPUB1EQjH1QWdrnoALwDXJ8/fOzAr0uwbZNSIGbF
vdv/rb1rXnHen1pNELh2R99pYX3LamTLYOYj2VYX1txg4DhAmMszxsMHSF/7AEU/eHxxZmLyD2+r
DIgHxp4UNwrNhNfYfhh057jUi6TgkxbCufeLX83WNYKa9JuezL4pd6PWFl0s7Jeu/ehbD+M/JFWb
epANH+cs7xvr7luezwXSvnYu7bnHuQCVjSt1Nq2FLj/uWUqvla36Qxc32vXUHALQsg/h4F2oT4Nn
ye7HRtR4EKbi+rJO0NUGoZY62D8mUw75MLW9qQ9hTXfr0SKM79VzfjcgyNh+4LL5xsy/8OfpwMyf
hpoiNx8XAXBGQYmp+kRGN0SiAbPtuSfE275/X4ZpRrcgimteYXrRE/6QcBcMek97m65XX0nYrEbk
szJVwqP/hUihfzonewYW/uDxHJXkyJxK84O2Dvfifyj6+uRgOCyO87Gx4jgLXxbKC8zdMqA0HTCU
VKqP2m73FFKpZ8g47e2Q9nV8Rwc1YTGZ3BASrVIjwV+ND90os/hfdhC3INVDrrXCEZvVoMLnzxqZ
gErtxF8XheR+54Q4M1juwVeKeHPjalWmgwJ3rtq/ZkIQPZ9BV18Wr9GKpbDi5Sbfm0FLfIPqMDih
aOw3k67G6cXiN4w16ohKQcDmwd0bQrDZGFm2V4zU6Hot7xYhx18ZUUmEHoXbHpkx/BtEqqxle+xW
/wi6jvozmrOCbIRGum3MplZt5BI0fcZgwtnXY5I7OGDZO01+bt4CcL+qGb4K0L6DzGhu7kg9H1Pf
JoYSBqEGXABXJdYQ8U04tVDuG8hWWZdKKvhz3ZLppl71LQhopncH9NMAJ8S5cNBOSO9LtCIvANEu
/s6vhMFuPY8BgAL3VFWCt7wEUljyUsCsK1s2yLhoUDBfzt8kW6QOtSl17C6ZlcN7oiu+Xr4QhQEs
t9ve0X/tFQ8jy3UYR6JX3M2fJRsRGmqhl+P5DCz1T1GpQaDU8Yje0FS3OwpbJS6grgHrAda0NRcd
FMUNkN4X6ojK1O7V6+a/dZLJG/+4kbaOCRkT/rzl9jzSaVXLAwsi83VZBsNGYqUrNNdfORCbNxIQ
9fOlOOBxy81VfDN1xV+7wx7rk2dRMudrmsygzTLBIhQSnykpPY/DS25brqwqoemmgeP0Oux9ghqR
USGhrAlLacYB/uU/mcMsYcQcZPBYPg7z7pn5RzzMrV6Ox/IXwI+HMTU1/cXRpQZ4k9RTt7UkxPuS
c4ukz+mOWdGyKb0ayqOXHTknVprkl2Ctqb4Lr7qcGm25+MYabCCElrX2Flehw4FbX19fmmRQ46rM
/ZHTKQfh9W+IHAcAb+jib9jGmcLtlUMy7R63QT2wKG4TNUHMEei0KDX2/++xnHSAFH8ebxFcQq95
/RrixZafpQ+heysPDAYLabJMPEvCBz9pZ9T6UuAOk7qf353rWPAn+g/beslrzpfwoWST4/GSfb6n
VVqxsvjZvO10XK8Etkr5CnZAtudxLft4KoeATAxsyG6atPjwU+uD3N9QvQOEMMP7uZWEzxH5mjGm
BdHlbj8O45dkX3F5YhRp0cqM5hqNXUo0EwHBax1FD/igCpnqDZxhkEm07r6GJQFz0NUTNKu9k6Vo
d2r4KkxBKPoxJ6Vkfv4m4MKD6LuRmpacPl/nW2zkK6t0JoQusQs8phsuEa42/9RM4qcrjSJrQobW
5Ha21sWK7Y4ahJVHda+FSurW0fhCvts73vV4Hev1pNUznkzAdFI76GMa3e9pSdZH6nfRigCDM1XT
TwdIgc3BcEwH083wdK0Brp1rVdQzG5DoH7v0x9AQ/FfsZEOW4oMu1mvKnJBTYUYJxUCSph6kw7Lu
HluI1+FlEVdFGKS99v0851+fKb4sVRTQAPA7BYRxNwlbQILmnONj3fCdiQmCsqRcc6mO4rr+p4iE
fLe+yK7gaYKbpbuNx4Fz1Tv8tIqzJMwXNDlOvWj0jIuS5I70ApYiDQba5uqHtL/875sZ437brpOA
J0WKLcpqPSBFa9rQ1bYwpfNlbSY1ZC/iC4L6tCB5eUUXAjKTtKE/AN0CyPtnkUUmvQ7gDrb1Sjqm
e/UOMHqgYO+9NUQJHdLpg76B9ur+l+/joB1YDW2tPa3dBiGoos1r9Q5/y9nkSPO24/g3QDYFkJMX
ElUTxFPRNWaAQP5xTmLus+fRCPa1iKVNm0p6pL7dMvSN3rnnzIhXHATEYLc/iACo0LphJu2a2FBG
lN9hfzWOJKO1B2d+7tTJwns6lyjJI2CwbgiQAN1n4OSIV2AC523nAJBIURXm1D77FagsvlMEl2po
WMgd/tTEYSYySLumA7i1JxrXzl/weeE1tQl31L9v13Xwg6QxOwIoDhb8vHfLzr/DTH9z2G7MuWZJ
2rmNMIFdKZPraIhpW3hEUaXfEKbSK+dZiW4J+0R0M8U1uaXMDQUYhvPNjOUjErSmWPNKT+qW+BJO
OsDxTTqK5SPov3tuI51kfVTJ8MAgLsk9GY5OO3oDsI+maRIp+M7Vng4znYvMS9QTVvU0HwyREJb/
VyS65MCXTuco/YibWGYC2Nqi/sgVXX/AcRL99WL9M6sEdATSjf0QD5nSB0a9jjDNGNOgEgzY9zhF
VpygaN4hg6rUnQWt655kzOAjOYFCTYgXv7YZ0AItW8L5S2EYeJwwqVhoB2YgtjG6J6BSIR+g2pBZ
qjhrThWEaGrucZma3jjxKhz7/ku9zdzOU77pZ8g6ekpbkNiCQ5ryx8nrFZOcHomU9O/ZkkQi4Gxq
VRfIqwQtEPsCyubo+Y3cRtTE2AEMQepF66qRb+I4n48qYNsEyvd0MBfyDJ5MmEt+EdcbBoaDc1BV
wglLtMVn6zpwFDzuqaxxXdn8CmlCPlx9GpcViZZBQHaBdRFAN6q5GiAZd4tejca/hQz5DAt4Njd5
ZxN0lw/9f/uggBLW3rzlrW5sDE5ul3W6BwwdcOWMqEsujw+cs67G8ilB1qEAc8O5ALaMTu5SNybZ
NukEWcFu+N5Uze/eICznGqx+/T8vtH2ixqTp23g6mabn5mfWN05G3Epw8TFO2Di9PYFOCZK3wGKh
agOR9+Wu3g2SLRZLXCl2QOjAvrpgQvez4atdAszg159hQ+fXwNbDmH2niTTpWB8wqvmHE7lUuevG
ZLeRajLN4HNXvQg2BtxZaHYXCDRlC/RuAsAwtl86PP1qZDqSV/ua58HiMAtY+Ah7T4/WdL8tfMfS
bcnCTHFDIEbw8l5g/aG4MDBT+oZsdy2waY9fWGHgQRGOYRyL/zW3bCtXjZjVWFNz4fXJYyT8hwrg
AGbSeUj9vs5xehzfWKogNUrdbfwVIRzopacjkLmt9s71oH7DnuTdCbMAaH2yw1MKpdarlyeey+UV
Wr2quzmibRvNI/87OIK31KS4f1Nq4lfkfBKBnkR81cpPdzd5Vo/FJWMFSYNJi059zyQ1uoPzEIXu
8Ca3ispeHm64bmVkNlnaV6T+L0MBQV0QAJo//MtyninBJ9whOLIFPqsSAwrMvw9+rncyytXT1Gzi
irBaDXsAwc/+L8eR36t1WKxysAzartyhHm8juhZVeUAXhH2HMAmAuOLpfmiTerq8mEDgq8DHPGYA
wrOH3b9eQzJ+dE88kgeAZtD2pJ/Q/xQPGgKtsp0HgsarxkplXM3WuK42aLbLpHM9G+oVj3g0wERw
Zhb+vK8WEqWs5Rl1Kg+8UFvxIdsWuSRtiVymh83zWPVr1+fiqc+JJLAvHZCue7hMDwdxp1d7RxCi
WCqC6441TjltewqAoRtT0aRC1nLxiBozI56m0tA7q3OTBc4xlBgTZ7X2P3VrhI45AsCkHaxCi5De
bgstLPpFIKAT3pwlyLxBSbLG59QqEqy6ov7VtfQ/l3TrHs7rvY7UxLnoI3pNJDGIPqJUHN8n8lXj
lSXXUWfzcWAo1wmTLEzumps+M+VA8dBeqlQXNW3OfvkRsvRbb4TC3ieuXt0gKMMIPlf65aszivSy
4tR+ML2CZpX0SaqAEHka9qFVPvg5PziC2qfC9tF0Xs9iDshBxauqQyWkxJvoBSpEgZQTG50uyGL0
Jxx3MnEoqa7lFujfv1nCTcfM8qhIf5AxUAo2cgdhVDNQWeozRGvp/omnWXGnNXBB6OrNTkZdPFmd
F8KDW2QrUG356BfF0s6Qr+C2zLs21bWfm+aDD+MXEL3vnBK40i01vn5Hlc3/jECP0x3YP7gdcfjV
M9YH1tU3GuuDD4iN3UrqaOUDxfHA8ks6W1SV4oGRfAHyUilkELS8crUwEmoeIxJ4hVDHGKOtW/Lp
9Hj2q+6VELXP4jF00sr7K/dxnpSKE6IUL8TKmbyJbBwTor5uK/3nz4LCltB5aVZ+LhQnhEnSfoSw
6yzFuAikIvaglutEMcg/vhJOihtls6QH9Ivy8hty30R2welaLrUsamrXRBKtRW4AjAv4u3EeKRpR
om2e9dbeiumirPpxDIe4YVHXZKbt/J8DKugCDLRi1I4wpkFiHf1JIpODHdMvOkg0ODjlOExV94Fq
03oJghojKtnlKB0eKE7vK1Fng6BEbu2uiI8DKmcmb0JLh390JLJR41BlHaDyuUT6OS63kFEIpczU
cWyfBALSfDzC/Sf1eWsTkIFar7w0v24+mfrv8QE6Bsaksv/RAZBUaFL2Wn+VJGewgNvqObQuXUan
ljlf1rePJmpEW7ppGcNKlrNu5/LzEt11+jNTKjFg3ntgh4rzDaE1RRq7gT7NTRU756MVNyreieX2
KA+gDGgdjp/inQxD75MVu5pWcB0lEaSmpg1C0HTwA/4q2ZhO5Cfon69EyZf46A2AYiZY/gykVhMK
6/eJ+qoH6b3qt350WYVFfsxyWv5vtg7JtscINVdBomn0zlHvtIxVzSxvHuMIobUEJhugt69TkJ/t
ZLBtnQ1BugQso+fy/Xf6EMyQG/4EuiYqH7dAuGJBfPd++7/3vYM2rtWmHwgAK5iKdL22ICkZYAqr
On9I+3DX7UI68l+nIbLoECNKRONClOAdzmBC19tR8miy5sUyiBhvhc6tX4Sb68Wx1CbjHljFItYn
/EZji/PANhHRsjllbLNsIeca3iCpErntdTH8LsJUl31StmJlxwJ/di/IaPiXOR/Emr1AyF2RbDQX
YQGi5cHcSntgVRyimk63vFdtfW8Qy9vL/grvOFR06qbfnE4AKi102clhdtuOOLmFze1K7dw11l4u
e8AXdQlLOr3vcesgnyLL7jNJYNg3aAQs57OsahIXssaWGo4Wx34BKBemgNruMhtIX53+SCKx6ygh
w09tPGlCVBBgxpUizg6lN7UkoiGWmgmRTM2tcbolBLR3SgVOWZlPjMa0Q4jVRQE95a8EOzvr3cW+
qxWwsJrjKZiak49FGDMsDNHjlNVdzXdPDjhUIuKeL5SOqv11HO4MqVFjbVaIiOcgPugF53a6ess3
nCgC8vg3dX5ihMiQynVe4iCTNaG4TwTjGq556JJUtSFPHxdwnjPxzzXdamFkJOs60l8uZKuZh6Zr
7XFtjCgy0p7OaH9V3mD+sTiDMmCZrwpY/GodY51uKX94OnOCRhWSrj5CyzyGVDmOrJqS7CmVl9hT
O5BcbbUb9mc6oViGaz1lW7gzYlx73tc5CrYGS0OG3l9EYsLpAHlHyu1C3naPit+6HRgsrxODsFul
zNR3SCI2lRSGy0pdJho8E5lDayksOjBQXvVlN+WaIM9Y7DJySO66vGzgHSRYmdVU05hA+7ag0yT7
FPP0lBC7l5aBJQZL4bWUNnQKc9HerihhNr2B4DJNVTOjoesClH4ep1+5bMy+HUfnYaexP2/ecoMd
/vsCMiKuxM3T/GUfgxSJBNPwHrbaBj0caw0ifgZthrBtl26oRVr8Yn+4SEF50tYIS0eW0raTDvUp
/aaCTmLNpsYgQgdmyfxASTFxW3RHxjOFH7PDKBqFUtPj/E+InMXjAymlI/CVT+8BOVZS00d/XB9U
tVFWupYyt2jjroKfVH6gJXttqukRcds+hPxt0IOnCLaOVj/MQf+a2IZXmjd8H55yJTsnHSC3BecO
It/rkVf+u4RXqNULXc7PmUEa/4IEcEp/Tn8BO5sGwbDOpbiHlxU64h9GJQ73XuMblnJRK5ovYV3W
Wu1/+jYwYSpcNDKirK2/Ki7DLNjLq1wHcMttrn+HNVWfKq3eZk8CKozvDrp+SCm/0bSeBSiSqcEA
REjNoyH/DqpY/bQhienBAAd6z+kwRwkpLijgnHipqF0Pts4NV/cEY5wWp8afeFjjJuPLxMrm1ekZ
bGGVp4Uo2A69crVKIQfXFdypA6zRI/FyejUZIST3Q6+EmVSXSGJAQ1P66slD6HXx92bfcL9Zrxkj
xaXG80NtzaGMImFeHm6msbniRaIRLG/QdMvGQHxozd2HhtSvGtXrQPFPEE5LJijFS2RhyYU+z1rt
1cnw37xxLnnyrHSAViJfPi15/fpGpOXq2A2+iHpqrjpSjpfuED6fgtWlNE8/Hmcmz43Tq2qGJbrC
L+oSAsSufIzHBTMA3awmeXdzdZNPA00b7+Vr7IXHuhXgbcXArmzM+eSEPqKgh+aw3k9kayDABosA
dAw9lmJV8GatgMD3/3tEL8Eo+zGo/tYN5P0L5I3dHbde1ardlWySj+KTntGpuEDs3efIXfdP3FLk
WntY3rzcbdJABezDQh3uX8FvpBQM9eKGTxOPBQZp+a7MhjAKl3y5Rp7Mwa2EK03QzHgtFrW93opa
cD8gZykF9NFw445vXYhpzYoSDXaErZc4pDGlZ6SDQiiad47rhfc4lRCc0DXt8aZ6QNitcPdYkbjs
emtUWOqWNeRCUCUoeBhK3SlGmEsjSzrGCpjHdZK5dhcWp89/Vicdwp1OUL5WOuBhaUJgqwEq8x7r
t+WBU4pvHmpNI2REb50EoKsv4rEgILDnnYAHkH8Nt71GUsyp7ogV2jQppnNE9X575ywk3Rd9lMdV
ASTNrVJgifyj/r4+gPT1fH5GjruhurKg1pE9S1+pBBImAyJNWBCSkzsT9Fq5ukT0Fj9O5ddlF869
V08HTkaVIF4wEVs+dwCo+7e+345lnH3nkTZpCV8571lWAE08nFbygQNOvq5fjSW8qM4e/+uWzZ+p
lIfJJBN7CsPEn9Z92XGZnZGlMH51ALhzsfN7pMayqrHoBwC0R032xd3iKNUYJiFGzshFCSzqywwO
0AWVGN8xfWXQnbnadcpfZ2xjkAxXTEAMtb0YJIZSFDb7QUrYXRTJmPzI6qB+y0ZW2n/oyMf6/ovG
0BZIhxwYZFLqubdlFfEc3GosMnz+6j8LOS7N66WNpP+V+w8l0zkPC0I9tbL/OfB7AnDPlNFy8Fwa
EYVOj9oBfvkZ5tz36ePpLUDWSOQEZT5mmBJrMeYI2XEZsgec1QSFw62Cp040eUIxdI0TavjD6LcI
mYjshf8l1gnJxsYCQyblqUg0Aky6P2WhHywIVrdGpRucUvhJqTbWB32LNfpchTIfQVhDUuBL7jiF
zF+wgSDGKxuBbepFFOnNTKKdIXo3riBD90fVftyfA1lYj0VDWt28hyATGEaEp82udlvm5Pn5hOMI
GxlogN/mKj2izJFihXKzBJhTXXZYtpwFkKkH6AwO0TZsNKgoSmqCBGirB+70mE5Q2GPVPmQro8y5
suQzp8QkaGij8bEt5DAR749q+ka1A8PZ+dOt+bsTGR4ts09cLUtKLxwDH9+NPu6kSfuhD06y93VU
AeD0RuhpLZAkgLWaAGSX3sON4C5wWAF4vYtsTnwcGpyLnHAbnofuubk4LY7iWU8ZDgqK2yIC9NLL
Uv8PLoOKY2vJV6Gb/X3VoOhJftLlFXMBl3GgtZzOQpVcC0w1LvaxFV9wlnKxNJHh5aIZl42a/BM4
gKLAM+K6YD4FWlRd656BTOLa6unWSPGznWdHEXKBrW2Cfx4V/pUL2nZT5rNlXSQ8Rtiz+UMlC9tV
8MZqTtleT07ui62gCpePN57xPa73Cl5vOXWiVFtGm2a22bINCDFF+GpQcY7Wv0h9lS+zMZOwUbGy
R2/6qlE4rM1ntN7lIjVjAMRwY/rei0/wHMkmYd7BqYQkTYHuMEPREOq+lMpv0rHWSGKu19yfwNur
iJrRsx6LvEIHOzSU+odtr6hNirE9ejnAuR2Wj5jVVcGzJal3Dnq9pHW0ByO990ZAf7492BctvprW
R4sCxB01HuykSYVoyAFAfvgAa/N0vh6cJzCoCpnnZSS5avLezXzgS58hP34X5z7Nck+YbD/jNkpJ
lYUhi3mRcTysPm37d0M0sTUZrU5tFk/V0rXtzv6edr1DunJfhEgNtV3kS5+JW1UtdKEWP0fd1Vea
l7Z5By6+6IPlPl9k1VgBwS3T1q3fOcHDxeUACbpVhnQhP0/abgL0cNHWXFXtd+VqKU59cu5y/mD6
WSxHWxcXPuiYKFTj5bvI7Q7O9usM7OmCRpYaZtFMNjI0bILYu5KSV3t0X7f0FsIpk7fUBow+oiMZ
GdfcQrKHNt2mi7VYRIBALVNwPxuJFWwNolCDy8ZZ5CaLCLhoMuCP79NfXNy1anrLkghG8CIuhF+7
eywAortD7kFtyqwYJiH/rq9V4pOZdHnV8FRJ4QZF2HTATSTksbi3Z4+79JV/yLcqcwWJUeAO/Nh9
4jaXg5rjdASn9gQ734A2m6/OdfcMMM7rmsWoT8ihCVFvbsnuOMJ4n325s6bgF3CSeFE5uKZLNa1V
ypxBtUKyr+6+5osknOZqgi+LxndVuIOu5MthB+u7H7gh26+leYO969Nu9E2UDW1P6FigtkFy3dOH
rPJ88DV0oXURviuGHHQcXPG2bPEqBxwugfpEu4psRxAAHM8H2UsexENnBYJ1C8P3qaNsi3wQMsDg
6arz2qQ8R2qGNQjJssDcH9cTNjZO2HEjs7u+ArDKjkU9mphcVcwZlbJxAKcseJzs/qwGnYFT7/+y
Cot/l1NfV7c4Fw7jS+z4OUQoNnO5YU2uFndQ0p8vbHADe+92l1KbushBUuI4ZVQE+sCr7xm0Ek7Y
aYx2ZhAL0Cp6Rf+iV4M2ODD94njVw9jJpc8OQJDTTvUpuePxMjGNqr2qFjnGEYRvlExBt5SzNpUw
wWT0t1OeoXSZFCZIRYAmtnhfRrUk3Om16SPtPDCq5bT4eXvxeuKK9UNns8GqM+7o0BEBEnbRJ7uh
Lilt3nP3BqpBcyDtIaG/XjaDHqqi6gQEviqiEv+FHV3ffvvG6eqplSrMVeI5Zy/nI3LWezmYeHO2
6tvrsB1VDwgTGe/nfI5xa8/dneyftww94+ap13TZLLcVrY+5Ol8T2c7Jb3znKGUA/RlI/oWiwBiC
GfvlU8IUvB301+nKjLtYkXaK9OwyKfs3/plZ3egct7F0TSxmF+OgkhHe3lYAtiOrSbc6BcXjEfUQ
05H77hZ9cBb7ndgAjfHIpcwYXnarosdfIMHUoc9pNyZEj8Zyo3AnEyclcMgUy7Weflm3ewha2G2O
sBsblbJWuqWjG46bO9RSO0nExCR3WEumQGQtTNMndVBwDBEdgwuTMMAo/uAm7G1I5m+wvCHu1E6F
xbDssu3DHCqhtJLLc500TJJZK/Du6n6PlvorD3NjmODVJdXjQL0G8cPbmWaFTsAFaOJQypkqZ0Re
nFBqP9BQr7cRLsCnbXLQ3Xv1YzSMs1n/ASNOA8ipgCItKrVPm804Jq5bR2yIQW282GFR0NCNYpth
dw/KdODwQZpi1u6HxLTvu6i8eFTgTYwus8Ru50Js13643TnuhGTkKCNHYAuk1INTfhlulNZjL2Gc
bPGIGMAa7IF55ah0mc9CWqUiANqrhZJyWAB2MsOgUH7CQNyx+ZI8OB2IRcBNG3aaJIzZLN1lhIP0
zVXtSSz8MemKCbVjTxyxUkOTuDgDiYMDL4zag6sSmeteBbkWFAFxmuX81mts3AokqP8SHbtR10p2
dt6Q8eQnKgkvabHZsxBIhJzj2XGNh3dZTLiA0T9dwMnrg84oJxPFoKSkccbX+KMpT0jzdsHC3+pl
09h+Yyzosq7s4eMVt0C1mbke+E27Zhk6WHY9XxiqW0+fxF7RdTn8z/EbWr2avk8/R/teEUOprII2
m3IG7XXy6jfRp2yc7JcDMn1NRiZcYEIsgMxKrQTn9xJFyJLuDqalUB/xGWqGGsJlfg3yUuJXTBGX
atXN5n7TH7X22esk30vs7FvdqpZExLSktw5MSdvzlej5qzK9Dv6/HlyQqXoDyljt0NGpAvp3LxTk
SIOfiztOPQpnWiT+dvO+ueIBnSQ5VslOElQ3BKrMDh10IHkalZvygHjwmReXhBX3wSUPMn7OUn5D
2DJMDtYXvRBF2ByIi5FyMJ81GhYkXKUia53YpUEz5hGB7zIBxRx1i5/emLo/+5hY9R7XCGozCuls
qrEIU/jhbW7ifw6FrtfTU90rRadfe5N0l1dQ3nd+l85HParuLoPCLoBdtOQG4Gl6qjIq5iHYkmhO
zQ2mNwj6w/BQS856ShO2W3KZGiOcDAjxvDrA/+DrfUus4kE/xdsFHP8xPcICIeBrHvweEIDwCtfi
bCIXvtKu60aDUi+Sgiz34JTSVOl8bmXsCNDEKC6y/bjQ33hayWi8IKK6g6vnIhw4F+5oW7IFFuFT
WenH7NZAQAjl3uJu3VXxjTgh7O1kBGelg/RuIpGFk1DH36R9w0C708mx7wEXGTVnng98khDv+7rZ
GI75MSDihoT6o2IGkeuUQ3O5a7BK+9nF+GLiLqLPVlVaZkGEfi4kgQ3dEkUR1X8104GbfF1onAhj
n2uvMnk7f/b/OtD6+kdBgyY6csm/nU1WzuoYo1dcTdCK44/fOY9nphhTiWsIllAeG3muLd1gk8Cl
VcsZ9Dwmr68XUpXtd2zALoV2zljDFOe8wPHSAwObufki92tzB7FoBsU1Cm/iqDKNMdMK4kr/8xF+
90mRmphyK0th0nfXHL5qjtkKC2H2ecPqcoT1kg6d9Tyv4riRk68sYgfXLa28PKcHYrim+DKj2Ygz
7BMaSozXVhTm13y0R8lekHW3qc2p8WYIG0KaKWYAUb6PzRyScinPjfnVmDIPOYKAkhz6doL/hRBE
51ixuY8ALW4yb23wGeZeFMFMEeZ/Lp4A7KyRfriQLkSt0N8JNbHT0vtI/jvbGlAaw3BvZBCWzPVC
2qiz4lk0hNPJ1Reu8kKxyusw6igX/XLFIfx73HHAalFc6l1KTRcBe3pdbAcMr9uFEwLoT4xgAB+Q
8cctsoscsCcxwKVYbOWUfXoQ1YUA+/B+uOARlP5xzWT2S6GVHve4lt6hDZ5OUl9/J7F7CE7So9Gs
+MPIm8HK5TbGq4tIros4AkGVn/ba3K2iIS13XVpP74ndZipISsWrtwcH75S9fYg7Z8ivPUPHE3r6
6Rx5IhdoK1EBJgO7ngSqg4cPwcmr54Fbbaz4XoKX3i/IYEC9G9EuZdL3ctl2a01NFGrQ+ILGiyZR
nIMi5by/jkxhP7kKfWtmCXcpYgeEUzivpAhBsX6H0pgCkRsHo32jD26Aokf8RMlinro8uJeNW08Q
locClOHIJAh/N8pzghzlizNzbuycWglXS+Lneox6S0f+yAslBZWbsrwBx+4Xeo69fCiiN1tB+fAw
TP0iTNkBBtnvVF9jjL8hg6In4w1EaOdFJmacfZcAO6CDDBDrxuw284pP5+Rk9eERVldm9Lp0QyWK
zaFoxJ/qN8frRgk1iyoPkD02XXrrjsHsCHEv0mJVWweeqdun1zyoS5iC/Mz5phNg69ys8CmgcJ6/
NZNJlEaYcRucj2wIw7QIaKVA+P+YY/rPAzpmCqP8dpw9fwJb8drq0gaAAT/zi3YK06tJDNamhKv4
wdrxFlqUJPYbcNg3JihHp7a6MPdEccx4bw8h+nl515byMPxxl/z43BVEj0tuaUH8aBum5i5qxLvU
jXR9NZJ+CScVxQce6fhbxL+GTtR4KZP5/Kvi3qP2dPwAwNxq83mHkXG60wLFPauzzFBptznEMNO4
NoN4XYVBQPOGU+HZDtLNop46K25P4WGAkUYYc72/dsYheKU5im8VZ0i92NbCEOGZ3EdBACLVyWKu
4Vq0zf/3JlfHM/ywi/gZ3ynV0C0FTgEO/g0Y3hIY2SPAo++0YEN6izSVhsTtxsvORIYMS0DLG+2Q
25Y3110YWAMaPR25ziJYOx64UKN1U5rH7n+xCjJ5t3t7hT8RdR1qI80AzbTIc66hsJj/xlCGltHN
lAyQ9f/VsQ35jjcpUTDsnD2ApobjUsB0U6O7xPpdOL+JAY34pwkLhxagEkzPR2oOreNkbsa3EsTE
VLO8qqYb+1OoKToKISXbr0PRyecWcpLr4YV7Q1OvFMWeozpwtno8mY2Fzthfh12okfs8EmhiTLNp
c+HzL4rMcoHWuHlpwjcrkM/Ok/AUOQVuefYLQLqaTPpMc4rERfUVWlDvYAoBXtbqUMGDzLj3afEj
zJ5vyHmSYSoZduJs4aooYt8KJuZbseukRntoJw3nZmpLS7olMlbRNSuOaIIMt1y8B9UphI8+jh8E
Ru0t9FlnD6sSTs65qGj/o0Su30TwvMjsYzl/axDYAIZ0dR8V3zfPZFQvUyVmCB+pdgGLOklOrBzR
W8IIiLtlCS1mZSydO5YROAP1yq5c2VxDw1fkevRsGIzOjFRnRsdY61bpPWiZJ2DUbm6yo38504RM
QHeWsJA8JldkvQhn8TWlK1j8basrn/Cqf2+ATLPYrxHdgf7p7EuhyzkP9IYsFOSPnI5oRDoXM+ya
Vj5ccPVll+gZd1N4wOljITZOjQcnpjj0Vter/uHCQA4fM5+HYx8IqOV7p5wLkF54mPn3dLqOZW8N
iyUkVX3bpZPlqYBF1laf9n3OGwLfbZHpb1pEIyWd7vJkoSbfw6+tQHj4SyEZ6KzbMnpVSN2R5qqg
/q/I3dIneBFxNICk0TM238bbR+OQgEfJwRm5ueHKWWMGuiUCqKj1AsT+bbPmAE8wXgskISrg6B9R
DoNTm3xI7zdUr4zdoMYrdITDyA7nX8+sVtxazifN5OYw0P9ZL+4Y2890eNFqbJp909EGpM9xQF2p
CNn1MPWFXTbKCACd7+Kh2SO0DTb1Lvqs2JDSILQnwf9fWrjZIwsYjLoVyXP9byK6wO+2ZR5OxWj5
wXTRaDCZ5ay1NMKJgE1CFcDXhahXLEwylqPxY67fuMPLYPUMLXom9Sd8FHJSZhlSODySNYHkzKMt
NijIb55+NJ++YmZrQjPsv68fjOo7QnqEZnsn6DACtT1rjhClhufwgRbFXnqf4VPWodKJ0tN4sL7N
uwYTM7hCv84i0RCxCyNf+q++mNI0f+mgURVmJGGPak0lWTML0WETjRHoBcVj8coS7oRXlYp3Ce9x
rHjMQqgVS4JL0ikMjKY2VMGen2RQFqzIsqd1Ff7vdve8mI9x0C1oJAc7ChT/Mvsd5LHsCq0Ap6gf
r6XA9RIBZGU0qGFIBN7hsGjIzhA9m8rctJe/u5PFxsM6FkXZ/wt8OrovWSYJ6yRejsziBUvxWjUU
dfYDyAFg9yBMYDhnu9E/m2iIPmzzbjIIUy0wybsKnrY3pKnKLl+SJGBL27tA6KTs2kuviFnX2BV5
/zMenFbpiePBXYB11yI145DivDw6BGJ8CA1bHZOatziHrgaMw4RYnQamZxY+8H7g2H19W4g/tKxp
eyxWEg/LbHhJTUWI66gp8IhPbE9VxGrV6ypFP9/bTTGt8gR1dhIXllJwVFl7Ust+pZS9MAFs+ldt
KiCDzRg4tKIkIOeGt9WJNOF5blXnNQiO8YSfvqRe8QInGBTXOtqFgMZu5KfAnjTwA42AnDnzxUPk
HZ3OBaMTz3GeXryPFqGy+Nt88foQhfZboEPVQNd1nwoWK9iinkQZUBuWYmqKDFN0BWSguKAMm64r
EEoVjwvk5myjjr171oV3iH7419+/ZD2meTR+HL8Z7z02rg1unnGssY7mplNHdl3SVc4Vq/xRNBl3
AkhqvsnW3goIi6TdebdXW9/iOORWClPFpfDj+ZO9B7RAw1egZ0A3DK30YaaTXPEGv0Xat8uFGbhV
855/jkpZf1b9tjNA3NNzPHr/O6yX3ftwlzAu5qogBpQa9uXEaGVWoqORPQ6dTE53//kgY3pXqRYU
0qf5K9FNQazhHrDASmxFWM/ox+yYcl4sNz9dJIyblqoZDcrIeh9DE0E0AdlCkrw4/KCElSQikC9k
5qw09WDYV/C0NcQX7Grui5uvqAVDDS0qiYlCTC0hvXR3ToZDam1Sig+1U+9OqvCTO9FHuclyJISZ
voimaemSmfnSAJ0fsqiB4vazJVL6LdXiwzBtLiFpcMEHs4rSBIfFnz+qRsyob6hMiGWfCYFUojtn
ISL6N2Fx0L8hEmqHtNwrK98gosUGbW0GuBiCh5aZJNfVE2iqmPttmHxNUXlccfnz88q8loTpQDAx
/oY8KA3iP6wHr2/N/6vv31gaJypn1O2PMqjwuEwKja5fcHIVfv2doXFO4AnAmvcgTbx+C1uDMe7i
J4eQYZ9nxunvnn87TCPTG9EtBkqd0jh2cmr7aFpjGtQak88cCSGs8abhte5ZRhJTAmrsaZjT3yzg
spACULUuJPH8HGvpx+LdgLAPOxsc7xKFZ4iEIA8by0ap/HGcloUyL9lW4S/eZuCX24EoSxl+ttc7
uhDEULc41ZuTOXya7FQCRpq5fuW3QtEjx/EITa7ZPltvxHgotuaAlU4/N2I3GcTKTY3bAnPg1eBR
zl4cRKO8wsgB131TC7/4XbFLlRRqWAusNqv2ppO3b8bIrsmuytTO447vOBpNuUWcMoh7Vv6ur51Z
ie4JwFnt/bmtZW28cjHdWA27qK9BGTHKFndb70cVrV55eetcHIP4BhpASUF2JHjXN307tCEMOY8/
HAuCDVVC8weDe9KshiTXwyP3RVHZ3TtLpXcr+TEINHXq0R7Zs7iQQIGHe6Kux30qGHq78j5Xzt38
rdjawwjHydDJc/Zkb2BBmXNH5RdzlD7VTARVfM5jSDcee785gl5mvU3VM8wnW5vbtg2ChcF4lm0W
drUFD32BAn6EgSP3eoEKCyX8Bbg9h7T5KAXFG8vPoy/tx8fIZT+7dpVkw82AagzqnwqY8Y7TISoc
t+l1vq4Kgrt6noJcF3PxTVUMAr9Ngb/Wv8o/KI8Z/pmjywKyXPqyJOGy4Ojk7p5neEgVV/Kaj8fi
KJFgW8sxrQXyxF7eGd3rBBWplidhnHSey2Rcx/y0t8b5mTZk6QDSJ2tTBBm9ug7kCAfXs0YeiWT9
acAt2QV7APW9QK+bGFAU67XzC2hDI1f507hH14Ut5g1MNbSOi2DAsbEo1XFV5aN7ntFrWnjzdntw
Ee+2mDTi+rXMNyiYQLVPHSQa/A7/5nFWlJk2zsbYa+vCcIWj27uNvah1+Wl9Sk9UX6nXT9VAsDIZ
cq0/48h3B1yZOvym5/IEv7BK2gbdxucK+sp0KlquA0ebnie0rhvKKGahn4qEEai94vt7rAb+sjn3
+3UixrNHSGiv7tPPr+f5oZzwVmKRovg8+pRFtf22e5FwgS9GGdoZnHHiSZaCRl0Jc6/mPAIZQipG
zRyk6UF8hJwpk71L/SUw3MfqWwwVl/J8+WVMR+wGxEJz+whpxWZE9G+8sZhIFNNDEF0KpQXCbGcx
hgrHc6gs9y/sdIbceK0FvkxUbLb2q3c9IBkDEZzNbibg9KyDacfmqgmUKIOpiII/kTyd5Ml0KLLS
g7AUGwtL8YsmGf+YzPRa/FVeUNVv3E6MI7NL2LmstGPVXEDYQSKI1Z2/L22QEb+DkBetRGJzlMVo
Dxt3OJY+ipPPcGPkYrg3JQz+m0KVKu8N2LqDGsef7Rne20O5bzs9Yn/33muEEEcvH2fFTisLjiVQ
yx2FFcZUEUvRkBRrsYeicb3+Llucf4MI0Q+1xEXSR/zT+tq3akWiA/xVhW/vaYxr4LTcOlHD6K0u
93mFJID6R/GyQECYvtg+qjYrQHdCjYccHv9zlY+AHJGHhKbiy7C0Kpxcawf/Oa/aH4gz4c0mpQZR
XOHJ2rTL3R05MfWSNW2db1wzFzDiMhTSF4zPDqVlpFGcUXsHl12t5zS6BiyUDRI+q6W+WCfwifsP
sK+IC8FIwfp2CWLbBFalIXDdJY3zV831p0nr1PiBFBHXsEKANWH+CWvs/gGVfZmBKqkoOMsztPKm
nhQwECuOgQCx3ck2x73+kQmlgkQR/N85C3cni0YfitfoKNlluQDmvqsfnz2yENk0fDF02lRo8O8H
SNKTxjqE8zxpmu4fgAzu+zWekChxd5MjP7pEQrMBPJ/64KXs93OZi5OAxi+VntrcwNHt5B4G9W4N
mq8ENQFFA9abGJKBMzF7wwvRrQnRc9pPc5vPqKSst2fjtz5/wljpfaC+zYuRG1+8MQs2Ov/V9/Vr
MhvLJvy6W6j+fJuTdvfnTf6cIkSo3u3cW3jEYeedUWvpkHQi7WsEh6dn1JOM7c5gKH5pcwudq5ar
6bSJ1XnAIVTQ9YgJLpImQ4jj5MPyyGbO9d35lHELTibGvICaEERyorIV9ZXJHPUMLYz4ihBmjwTc
q3iAt83D3wWCxpf68Q79thKXcA0Oml0k8RIglYhxWuDdo+29u+k1EbZGmGnbDCwriXoUbu06u+iu
gmKidIlY9c7x9W2GcrG35Hw9727pHJ+5Bkvzx/MR56DsRY0/27zI6ackvzDMNBpH0fVOpKOhLV0T
KKcQFMzE0l0PkEVepAAGehbWx5igXE0seiJEHRk/FA/cr/CNZREzxxxQ6tGW5JGV+lFGjXGxgNzM
cEQWW5B7AsP/ro89zGDT80n68DJbSCGcp9F2XwH4RVgGjCPVPOUj2KtNQfn0iHEhqSeOSrUS6E5l
666JsOgjCVRiQ4EQa6qdvIzR2lFxNgd817yhGUu4NoI0y5fzKkhCA5eVQNHYaEyA9Hvo9wKVYNGH
MkjQidasFZpChb5kAJjJaiJmTLus3ndGCuWen+C7c2CSRa+zWIL3q2CTsOL8JfYO7iTOpC1wtn2K
YZGodwpx8qD8ZWFVVM/+yxvQFkzjmkmNrJDT/cIaBzdSqmwqoTVqk2UNI+NozCz9y8PbyG43kMO3
zivX0gDWMUNgI/Bhq1cS62BO7wvc2oBQIqGf1xKR/rh13RwkkIQzfuC06qaeikxFukS9Hl0EhLuh
QwhKKP8mBrEACNPHgGdvXm6aFJN0PhpY101FwjekVAvppHIWEa/dweC35DcieBZCtJB8Xobcl+UI
mAZkZSMXuaWHSjJRHPydkmFhE1jVPQPnBYTbBoGmvvz3ogpHE0azz8+ACk+FkYmjwmr6L+z0AjPg
C8P7bYZKO0aRPw+JN5mB6/tSLyx3GoYxhOuPcg+L1IxGJF6UPu04JiVoRy6+nD9f/iZ7dmo8JTAm
xMz2487+64hBPLxByz+FwlgBf5LeMLkSja9UKup/VnCSG4FCC71NWxJgy9HqaWg2kBvIKnqgwg79
zZf08fFmpYoOLg28ks8JIyOMA2N4M8e4/gDpDDJpvF5JrVlFM6Ku6c65rH9z5kX0I0ZrGDyztQnK
NQBFrQRT41gdLHLTj8grYrAfihsSoYjV6c4ZIcFyMHa/l4+3A6exCyi15ZiBVNJFlXt1gOma5I7J
Yq8uph2xFIOf5AwT7g8yQZHdXwerPs9tZuuGHF8LujJq6+4npOmRsWlTlro0XYrc2t85agXuJVLT
A+hJn8KRkdvHA94IiMvDLjvtR8rEkWC8dmNwuIty0OS0m3F24JQycyTN8B/2HG0ekv/9NtOngJGn
IR4J/XnTh2C5aQZUsPYtDm225aP6IySOV9IEaIojHR2ASlA2Zk1UMvoI2tdZ2caFpMsgE4HaZhOF
EmEMLVF/mAd4trNyrZ+8lYwTPhkPDtE/udnEe4jgtrkWSMa4cYBngN/jG6hVEzSHgb/FwrwRLy3q
WVmgcJq+oC0tFS/J8jaH58X57NXoRSDSV2aMRxAIezxLKTzgCBZFoR44NoGyurtAl12v674vgBWA
DVZpWH1j9kis15tgxi/EK0iQgim1RR1tY+0Dgqrv0W4mZT4jl8lvH8YPyGHxfN/T0LOlgaBbDbf5
luayqNdhAL3oz3nA+xj9ygfZiLjZMKD+WcMVS7wAC6T+QOr/KbszIxYQ1xpwVS7wDm9zdSDnGBFU
OHZrSqBS2mwrW3Rd5G4i4DyR/EbBd1D9MfvGM8vRL72SQSVsrQ9zDGuq7lGC86BQOxc1hcR28YN1
Te9tX8Mjd7pKXpNor9u4KlMvii4a5ZMxiNnNas0ks34c8olUGAoQbvclm3K4JbmYqT/5ym2FTyW3
KKdDQWPWhyCo5MnqU4E4zb2c8VmTvnrvlzHyHgJ7+RbOrNY6ddXQHkkdrOOdy4mcdMRF/fFdG3hY
ZdZljKGBMlcd6bbUIkB0spbIxGxCnxpGPeVv4G3/6FsM8DgVnwWj3C5VzGDWqB8SXbd+OtVt/jst
RH8LRdSnAw52lkaQa53kJBmRouWVGsrib5OCEeAIdPHLRbbGDXNODE/m5/kXd3x0rLUhsjxy5Fch
1qiuSk2Y/lyNEAlteI4T25HoHQUzg5AJKuEhkeIht3ABrTiSXn5dE9PQsjxl236/j/tk7VH6wbfp
hfPX24QMKErg1nkZrAoYCQguck6EU+Sr97yqSsg770TX6DeLS1p+yXF4KNleb2M9M66bFUJmaVpE
qwj+QoR4vQMxV5eRleciDfsUMw58ilaWP3ZKh3e2vr0FDE5NOFz/JHzMVyAPKt1/3k1I6X1RzI+/
Z26kUuPirTUPFlCP2ONZzEBrmpObL2U2lyK8Or0qqzwDOO1w7m5J39J1EsMWLSzeonccXT6IdL+r
EOyagVY6KCgO69ZvVFqK4nv22g6mdd6RMNoJxIIea4/R+w0kz4puqwZlacJVtMpyjX9Bd9vR3C0/
o09lF0hvmEpOk2yEpCzhINHMXWnXKU/TH3ehE6Enm2IVowqcWTD3so+SQxv27IFkkwqVuRMBM3ou
cP/nPQqo0FYgku4bzeFcW2/kdx2yaePZVUtH868azwLY8tiTpUyzw2PiE01J5xusX6v5GR/nLlUT
pp0O3o2rlUYg3RlBotdmf+ZK/+2gOyqu7VLWta/wXrmjKzU7q8qlMJyEIQieN4f3XEL/i6o+2qmN
lM2XmzKwY7447dJljrQOTKeuYOhh+fZV16LXpIrB4faK8Gz45acyNq2a5FC9FvdaOMKBI/7cGOoi
2C2FFBEZm0wBqxUvujkGAjD69S1MDGmpkZc7e8KuC8qhYhx97l4C1Gmdnity48UXfj7aAbxXdUP/
tItv1321NZnSZ3B7pv2iFvq5LZ458xhFZ5bz+EmnyytjzWD9P8wFTnB+HAhLMtbLybIMO+1yUQpN
99UTe4HbiNIXibNLZyzGUpRKf6fCEWohTAay4e4bm4tNtXMxY7fEZxVKAJpjBVfN3lAdLLA305Eq
+r8Oaqp41NiCZ7gey9nKOdVVboEd4hzqhsRWkhqSiAEwViZaSyatu8UKtQzrQ/V1J/tIFUKT+tLC
7+dfXWlVufD+ykHIXksNIB4gCpjnGwRV33Yx2nli50+rFlPjC7kOczjJXoB+JrX1GwV/usqSNLIJ
oggJ9KqR6uJl2Y7vERhwNPPrMUL9NJZHBKrrW4bqeJGfSYIeMgsPE9LEqAdLbqcH86+yZ1yRjkGR
qRn6M4CnaxUUp80Vqaz71JAF5wPKqPxJXpcCLQW+mb2kN85E30lEs9ZyUZawmyhI01ZEKpsnZvrF
ejs/BllzJhyfoVhdzHP1QKEZtyof7l51uXwANPyE/25HywU01sXphGXhBARCQfdWKEgh9NGSzjQk
+81fX71s6yQgs4ZJqHzgn61dnYbR7JZJojK9VRFi64eWhiGklyHN1UXKVQBgGWHFTnU6RGWwA9x2
HBWuSXERouqZ+pb7xMuBs+LUJ+kOH2pFfM5NkOmzQxw2r+8HVJ9Ew7jdow0QL1HkCZAPNDCwetp/
C3YI3XgmU/qoL4C9eZdJ2w4gRzJvqV0H+ZjlcGNxIRs33Abgpt0fQs+VJE08DE18DndRV7i5Rbgx
KfelWvGPh/vzO7CMYZ1KW8jEGZnQ3GgLfNY6kKH+tAOAF3+hkmMUIURiFAu3JWnYFgCok/FwdXr+
3FaQrVY+X0cwWjrcNZhuD9LCnThgXSYIoFaENBtQwKu4PI/r6GwZDXO8kii8xu56sQP9UfOAuHfc
F7gO+UR7iHs8MKdRB0sCZHBmgFOzH9UceJlfR/7DKTCshGqOkRw4nPzFsOnFfjQ8A//amALY6xER
PtLuZcuIsjE3C3S5lUzIkPu2bXYUzGOMpDdAb1y80JS/PY+848L/YT71JAPYJn3zVQn4mMPZpDO2
tteAZoOVpRYkQEsKA2rHt6Y2B/xM5zQC5nTKL8HjTdJK7SiZhu+nF2ii2Uu6OQrZy8wKTZBjx26G
o5tU6maUEsLuoWyt0plYvc6LAbz337rHOQqaL1k1bdHYt7ERc0VAA/r4bxEWXh3z1WmWa4xpCho0
g416XqrCZ4lUXaDN2XBPfywKbYJcHtEEPGlYwcwN7ZgmvfCB0lup+ySabYQ0WkbNGcfvUghaPZxO
1gpyoz6vAAr2IVmBvCEaEzVms81Rf8meCvlZLgdmoNYYEC2iayRNrTMCjdWSCtP/7h2sOoBTV64X
qay93Y+VIFuzOGL26ZO+YgAw/eoorwn2iTA4Yu75E12sPrGCVW9YUNIq0kOBZCS7I+YVfx8BVLA3
FaC4wMHgS79WhC/E4l511fEd2PycLISJ5Vw2lhLmX0iUbIv1nOZc0XO63gxTGYN9X4V0NnTtyaY4
8cIZs3jEi7w/2G4oXaQenoa0ABaj2mW28zGH83EWAawtjTqGCoiLSgJ/yBN47ZCRtaCtYyRr4JPA
4cwExczTxC+G3hfgc4CP5sGFgfONB7zJih/P4qFrzCKocqmDMWYi49vlymnkluGfurMXXL1gyPUs
tgzMjUD+UmKuN2J1FqyMx63UXQrZjs6IkAZZBP+r4rWAdaF1eKgoEfR3dBQrQHYg07wdtMdst41j
ZSTddqw/F7jUYqEVx284+8vAhtEg4dS8dA/M0SAEeCfeu9KjQsyERr6mZwUxkgGC4ttThKppfD8R
NM9hZGuOGjAw+Sx/eVwq4PJi9W52/hi3wUUzdGmzag5wCji7huHBhIxTL1ERO1OSd+khwfHXL8fz
Kwjddtd5pjypXa5mylbxCCDQWGrOIvVUmMm1pUqu9R8I0V3gkmmLJO61gg+JUSxUjxRPusLSK536
ZUZmHJVzPVPzylnpIZ9td/D7DN6hgOjWDXfl5UTdIVaym0CSaD/H1/p/q8Qw/SnqduK0P0EPG+M6
fF7+pRmBj5YO4ph3aGVaOwvNB7ETsRoNZbnJkZ0W1zrRfGXpQU1ZCzG9NbipbiW8mHv5NuwYmJZr
bCoaap8OE3anr7U2vr8k2JWtRm4n6Fo3HsN1GbmajISG2mjYuE1yM+W9QEoR2gA7YeoWqr+fa/8A
3Jw5tww1EeqP7SbM5hq0yNAPhFkYEDUAi2oFCST7l9bj68Q3eP5Cyj2+Wwc+SDMxl+4C2OGs0o6h
ujMZ6g8rixNIsV9Oh2lSMk+ZlSvMtLlbM2wldovsUtijYS6dTmP3AJRbtcbPTkj2Jv+q8dBcC5u+
XTcAe18FUTrhxaM3kpEYMyeohQJiI8vbcbxSh3YMCiUTcXexwshiMYbOjIGzGsHJ2ojuhkxduj56
xNDKIIuJxovhcskg0UNxlhU7eBxoCeB4CSnR2BmqWvnzmIwHd3yHfG6bH6yWRiTriF7VpLvue2j6
l5wxp7buL9hyPVAtS1X0Ef9H5eyMww2F3kljVicuTCX4mvUTo36fUjlPudrEOFOj60aRNptmbTp4
527Bvz4+OShRF5m99j8oeh6XUbjGw2ewTTRniZDCY7TQTeGofTc+HojfhFXjHVXKgk4uMeAJHjez
EPLKLnWJnzRsD+hKdWw5gmNC4zXB4wb0l26bJzKjDjDF9KO0KVavmAAmNQh2HBTkhnKTnyZcVJG9
sQb3bZoL+4dXGH+MpR8nBoiuIxZBIFzBkElmV+bWnZGOznBE3lfNHeNMcAF2jtYTXDL6hKlIy6sG
mb+pFDDmLNicAl0PjxJvbhjySxJ2ZGPcrqfcqqTFrmwYSA+P931bwFE0W+/Z7UWBvN7dH1p64bsH
19clPL0xkxrBMNSKmjuYxvjkYCBW0133+pnhGadSNjQZ0JvsLXocTCl84Jt4B/GG5RcLQtQLanKW
wwoAEGBhjteTofPpBCoPXI95/zYlitfecJHF/D2sCK/0wPoBr6cIFGVyAjBHkMYzpTa32QLqs7vK
6dDh2ZAyAUeUpsx21A1/9m8ze7tbc0G4CylZdWDcjYXBsyQKYh1U+1q1bGrmYmL+LrB5EBZXDPOO
gsHhE56Csil08Yo71spbUH+kDhlcSDYXdhsGDQyM+QgW49McUf2WE+WzzM9UELOLBd55cNQkX4aV
FAnI2Ku6ggMJ1P0KiJJCZ6D/5qmG1KGc3aRMXWs46NrUUdigSJucgviIMgXwviiXOu8qcQlg5iAY
lhQ84zAH/MxrGol/nQrg9ZXmjBvr1Kooog2wDtqWntB1bPyo6ME06C5NFCpT9sNuBIPu5HrK9hxC
l7ty3f1JDDq693WxVr1JbBNGQRPpBQMmNJb24Y+QDwNrH2lGzCQyLcJCSFxovO2+8X1DqdAKwhjJ
sgnEEja5LikOMP0eHkzFWTAs+VigqPx+sFY5fWNynDGLftQgTjVb6VB2M5A3kxrL0SwVUqpXYEbC
AutY8LDyYpvNKuOCTcN773r39O/e0Fd0z7r8yyxXxsvDiigcfhhO4GhIcbdeHT97NwbrVcJ73BpL
zrNeeRrdAIzNtMa7XqOyfgSDF/87vbkKNHrWm/tPgTS4dg+y7eDu78ciY8Fp7wKdQgC0zJJ6dBxR
2RpePy1ulIXFK5S/49saIsOZRI/XMwngp2iCaNRg6XFf8qT6/4KaWG2SCjmN1v8EP5fEz9BkJ3ye
eQnnEp23anBMGRR/rrbOYROBrD1ae8ZBmvg/Vs2LpUm8SK9cbGwCBnvpPAOLyrfNSBxcauf8P5n4
WuZR5OYT2bNRk99wq4biDYEOIfRUc2CTxkBwoAwmbUZPPQKcn1bkWHEg3heb4RctrZO2TMUjesw3
JYJS2CSoUYqbx+XjKG/wah6HiR7dTDe0fRtIqg8wCbG5fFf3+ObPiJcEOKKfLyvlSVKCFjJ5jx58
CJTvzNu2kP/TOcJILnjkQlqg1GehLB/FOjPGc+EGZbafQUXTi7fp7tkyu7DZmAT3aYHFVK9SEvSM
TD3chZYvMUPt1vXj6JflaEzIXXXkLBgwBDfK2iD9OHhuiKL34U9x8EG3IbRHonq38xwxZbjT5/M+
sd9sh8F4IcsXw7yE+gBp2pl8pkXzGxUTR3UzyHNcAU+Ea1jxffMSTW32oZXPbzd/pcrA1vRm2wqi
uWUHuOO7EpIrw7XZ2dZJl4JE1rpjNjTLtGed1/dBZjuiEcBQKqT58CoATwYERqiADtT6EKOIph33
sO0bAZKp4KMDsp7hDW8NQKyEt5/XgPwf3N5C1WzJfZ3cp4CKZsjmlWAlgf1RLMu0iNHxlEeo9Cax
mzWLMld7WCNMfYT2dfP4QcOPEIj0ehD/ia4pzgDA0afQU8ZMQcCKrHjbtePZKO8hwRVS7xDE7yrG
1CBqFqGjvDCd2+vW7pZmby91I3sBW0bgMGoq0sNb+JlXweQvy8M+Nz3PQdysDepitKIgn8Fc4nfy
6WwlBpMO7QyMk2AlalWnRH8PUSnUAVc6JkIHUuqW8fRdVabijc+YQLcoPRUMFuJ5YVusCAlsHKjY
ZGaGkCZqZJOgJzzQlzxX+SBiF+MOSqxS3BDtG8IjImxqwNxZW299OqcadH09LYqlUk0+4kli8Gz+
ud2rbn+GFrO5zcbpBftCnXDefaH+gu1JSMfPGvPU+Naqtj0hfcSBLH8OevEzTvOep9Y/8/mRAfPn
V6WsPu5ZSY65W8c8GRQSEpdwdIjnTRjWivuC0HspbQOw2X7HX6enPE7nIbtsavtrNETtspawT1C+
KpJs1sAkL2Hlk5qM7hPuHLM0xLTJY97tXgi9cUD+5vyC0Q6ajYPO9rvZHuF67hhxMpS9e+82QThK
xX3OeDGLrAvkGqRugvzcnYdNSwzFRF1rvTstaoAeWzaWisRSX8wz80+NjcYyzCnArpqqnVBK/79m
x1L6ZsAgjpVyGLwWbxetweLtiAKVtjZByFsvhzCwqbFkbyHY1wotlASXr3YYTX+hKE3bRm7gGEPZ
eDFP4RqnXx6czfHIjGfejGXDUkBkHSSkr3pr5/2+UPcAUQOHG7tE5VF4TvCxqKXonmTVZXr8gox9
6oASvJzAkLneMikt+ctRC3gcPhh4He20nVuG9ihwkrGvI6Zn9A5x68dSX8KCTbVjXgCOBkFIWvUJ
JlEBe6xnO/mdU+HSvlc2fDiViymmz4RqhG53W8s2WUlcOBGYljxh0MqrYVVZqYujmPFaQCOL6jDU
L+9K4FkR5TjmJilDxVJk7yxdvaIdTaLfWRuNJ/lzviuqWpyzrfxC6sUqMw4fjuVgCHA3/QGV0Jqy
9bCbfh/Wx41yt1JZCOoppvaoVAefZNcqJp/UaKZ6Gsnw9oCNHYD+socw4jaUkfMsoCYcqMMXuLdB
8/G2u+MOS7xfGjPtzmRXyofU66y6LQSnhzFVjRMEmCjTKWB6uA3KYGnigTJhmxV0hhaa1FvcMNdX
92ic/j95po6MDNQCGKK9JrNNSCQzWjIFckYPKEcixDzejH9JeaptdAlDnjNnB/bEZrHVDhp5iy1Z
AMHlQjy2Jcm1di07dwEkVy/0zjKjdoQ30LP5fphHFm4UxZ1+0iY5qbZw3+R5DQ83axyLjuWDVYB/
0xrU0sznGr6tPpeGQ9dxQ/uSDhqSt2LS33fZ88DIR1tCorz9fDjfOtlBZfDeDI3QgZ6AF5Mu+a7u
qS2EVWxSQEr7kA4zNAf5A4RmWRlZISFEtKOaPIXPjWwLsNQMaDEYIvsKbNiprI5LEK3Gh7BiCUil
01+tPDdYYgFjiTaHnA3ViqqG3ePVf+FmHdBPSmorO3yDJB03doLrNWfhHFqbOjagGW9NpvcBsNQp
wo32bXoMSYD3Xxp6lM8+29VL4q07F9ciWSBxPuog9kKjnXKoziVE8kKImWMlcC9DrXXdAb9qdFPK
+9BkARbUYgEFhSPaB2iWk9cCQqLy1ymG9so6f33+jTTBD8HPn2y4Oi7q/AYlv4WmB9TGgAbYMGv4
mWQPCpte225hZRWkN8GPDjkq5uAkkM6CIXzJ1aFq68PQAncJzdAvjjOU2zqgPBOWjewMcdMje+Ix
pqyx9SnuYuIrRXWFSD5Hl//l204SmKrsOnqOqTiAdsAFoib+aeJ77798B8pOOqZI9qsI39rFNsw+
Iuta8y5M5kABuSHOLOB5yq9R82IGT4V5egoeXGDotCvo4TxPwkZnDRFxYCxRRubpd7IPkBe5v6ej
Nk36c2mpbYr6jxCa9UUZiyUHlnALytK9QbYQtkdaIsvQz9ta/iLvCy757mS40xi0DUE6nYJuQu0o
XlwVeTbqBV0/mWUvs2dWKaDUHajQ1FkNPGj1x3AuUaedKS/om8bd7w5boPYNe04NYJDuverE1n5g
dHFY7PCRtVJy9tC3Sb7vJxDR3uyppd0TDIc31fpH+gJbAokoK5BLX2WjzOSooHEe0qo5kS2E8dt5
3kI6XSsDbjychyy5/BjwJEUvpun9izrU4EjVH7MssEWUZ4MfePIz4+6PH3e8otjXQGErbcqBn1bZ
BvwWlUspNIZjgdrTwetE1c6qe4qZoj4UNZ0N1q8L/N/VXNoTSaBla+WtfBbGuCHGzTbP+fOIIiFu
1Whltinntnj/u0puKrKIMlFmdIMAu5X8EfIDCLV35VqjTqPbQSfZvtLkBTlZkO7PPbjwFdX4KVvp
DxuJhGdxuoYEdsO27JZDyzb3LWTJbd9hzTu6Rs5vhdpYtSebUAEnyJ847g9Q4I91tDvLb+JukALU
jSP9DTgpsTS96M2wwyxxH0neJRWZ2vEUx7blKz5Nyb8VtpQE2i66rEyM4OJSBck08E1tOhnzEzED
Bnz5264Y+zi4JEfLjJXrdDgYo5LtkkUv5hDZHWxC2aN4mj3JTepSzrkUQ+sWgX8UGQ0anoIdOHI9
TQxOzQ+eMDApSAxb5v8igNBpx0slaw3tDdleX7HMTCqicczxOeaV9dg+M1cJJ/V5HGEHBMzNu9bP
eGlmM4Ci2hQ/EgnjTgtNRK5RpMX35oJnRSVKmxunhrKfJr5J1GL68Bqv+2U1eqfDi/R4TpGn0r63
mzIy5Dn54UWjb1AzhKK9AcsXULXMQnqvlsDSX5BNLrJLnx2JjujivurDaHdv8YTanPN9OpDcyhzY
bmSeDaW5cfXuthZWIJm+lfz5bsZDoNGWyYMtTbvwip8n8EJK1JiaP9L2gDlrXoiRzgC2GeCrPXDi
aNIGe22X8R9CCzFY9so23I6WAfC0I0hz3Dz+t0gFLWt7UXUseT0lQq6HHUsRMR6Bz1LjdECFYuOa
rh3/MoEOKywZ1rb5Wks776haEMVW6fTg2pxvkIwIKWJS85uM3eW5A5LY++8SeHEuU661Bl4rQYfi
A0gjnO3UsaGvaVEVqL1CHa4gJ3mqH1ivKlplKwIjO9B7IEjUOHEStuxVqeWTs8NMU0cjQW9W+LdG
DZ9hQZSMzv60rKzWLlD44iavYBuoHsq8vluy1S/OWBIWI5xGfSQtuPULN9Aoyx9oygiYGjbd3fAj
Y0c2n3iGOL4xgEYis3FVki7Oo1YqQUaqlXTiH6I4K1zOvUfQQ/mdvCBcDzlmmCDxAPJgSt/0sXqX
CQGbKJRE9dABrEEMaSDb1yLkC2uwsgy3kcxkn4lZDvDXKJ0PH7dIAGwlGC3JJH9teAoUlQMlBFhd
Ea+YklrPRyLmjoo7U3Nz4Rm06S8EVKUviJw8kxyHpXXISIX/NtHMbNSH9ygNBpyV9AZZN4Fv+YLM
bQ3/bjatuNbdifXgKG9rBY9v/bPJXXIuQalVCZ1cOpyox3yumt1yZZOtAG1NxUDuiPgipYYYmrYd
lu4+q0S/MP0i20Btj6yO/7xflVWcd+CKsLObQKXGxELZX4A+nmHQSuAom+VoXr8OG0gcbEdbsbKe
d0zIfbasdo/LrWLzc4w0dpDkok7n/C80Di2QAZMmGTuHvmO0ZsBYp0Uwn7Rg+my1kDO8z3udtcqQ
KzNBxrjqtMPcPy7sX1RCbTkQJvults85oQg3/ry6Kcu60EwD/skzO/fD9iWWvQf7PTdaobLwsG+D
Kx3T1R22hNfv6s9low2Ovv8U+u+C+EWfQwpE0dK7FimkblnYdxRKqpPsr+nrFUr6m1e5I9jSUDDQ
aztlXWNk6f+7LHfABRgbiE+2WRR7F1ij1XeB4rwrWmUw6UiLeKrQsibKS51c+9C3XxyjGBjNUPx+
skdllru1ktkULczUW0yMDYS4luzWk6oS/8Mu+SH0Nmcxrwew6QNRjKXHqqT6SXEluLiAP4lo0Vnf
3y0zfQjET0yJW1D6qDUrZgbv/KvC/Dsp3rwZDH6g+D0q6XqWbPR8FVsRM4v2tEcwtyBjHXKl5073
CFZqBUjRnZVNXHMdji9S3lVT1Ht1mg+nLyMWkIQ0Ew/7GhV6eMDVuaLw1jT0KKJMAHWf+z6qA3E5
wcUQ6GTErXuoUrQPRp+6AHBDMf4KQRxk3i+cQzAT2nHjm4RhTpooh5k5i8lKkIzQP/demcVBRAZ0
xvBCLDXmHrlBjIUygF5gnRrjgQV8ueKULaumd+qii79vTaN6r1yMf6A8kLVTvW44vSm9kTWp3aWZ
M+tpoJtiHdlBCs/I9/NBhEEBukpl8cXg5y3NoHCUmJoLVR+PU+r07wbP8KszR9Agx/y/89KnNewM
WTFjQvSiIypJjHIswuSMuGZcymfk/g947EqRuln6EFIlsq3S8GlzGvazFZtEv77lmXK5zzh8XJ+J
rKB/loK5IzDIjSshEqfnEO6nmirKDw145XWoWrqHoNCpD2LgLelEgJnk8qTy7OOl7x6EixPep+y6
edAxT0rfYeRpC+a3nv6XgIS5v6kqSn3aHNeLBrG5mx1mpHTYVHprzqUQ2Nqxif8Jy7IHqNVvay6U
hdlpqZa30QCYkUF/BLnzY6/rFbW6DmlXpa4GTAPsMxEed5xP/rUMRjFfdExwynczk/A+On6KF6lq
nIe2xqmWkrUpkZL87JdyTSTy2wpY7XG5t38UvfKD59T3Y4EpmeO44LFhVd0AAj7qgQcGqU3fsrsh
92Pvwzw4khYpjjBX3/PkAWJHJlp9OfsU5RhPjAAtD6UWuu4YDpZCKdMnYE9i90KBRUh8GC2hbQ76
VmsZGUhs7dWwUAie4o7i8qyNPqK3ZhsgMqIO/cILAcpHXGgmTzonp+ml5AmUILigP7waF/GCprAx
Lc2XmXEo9fBkfWuA/48mkCD0Ds4vQOMeAABRjatX9txh/NRzWMaiD1AG4i/ZoSErClCie4nAJemH
I8eRljXL+7SHlaSxVUfmUo0WzI9D3g8bF+EZjegYW5h5lcBaLwawbbtVv7ao1wslxkYyjExIrqjz
QaZ9N8ULs6hAV25yqKferAEgYmPxypvE7ndWU4fUvUVXIWptJaaWy18Z6Sx6FnNDfU0xH84u1V/0
WGFFonKB/bnV6Js/akmUDHo0kbNnXTF3qXem+N07zLPdc+cI/yB9/VaDe3lr2Q66ok22QiImANzt
L8VmYHsqOHkpQtSaoaKUJfwbz0xUAxTprXMignWE2BxyBax5zJC0kcU4FC0bsXFwluBvFV6ggWsH
32l16ngQYSQMC8egFu0Vkf2zlLPP2f6VDSOjyzoII1jEUP5Oh77dxrsSGvGLJ0pqWshFSPy2vvZj
TXJtZaaUQ9opozFHFtc8iMxJ8Tb+0TRMaP1alf+n2Gu8dxcGOcbYgR8EHdxSMaFS8MQ9Hml1tM+A
4uvBOIqtaunvYRUKcY5T6kyS55ydizWqbOP8WUzxC9Fz6FpEtKcKBXu65gIhRqNxrKNhrkGwnAEv
hZyeNsZFeSVr4UYfsoJGV0wUJCO9t7YJ/eThlj1P/nBONFfsDljLrS56PTHLAwAMCfGGvwUxWv26
P313brhKNcKPTKMCernu4QGfQ7WsQtZ8kVvmzdiaCAftQ/rUceO8xicOoJdPPYa15mLQ1obJ7H0f
St2+Rv3r3ai6XyFaS3L9xYadTV5NjJaZdQHvbSKCTLbCDp+MhgGlJ5AiGLBFiEzZUHeAJSEOWhtq
KXnaab1KTDq1YI/pugr+iSpQ0gL4gjJau60NArH3ShrPOwoCKuPiKgVxZJ4uBS4J1d6iPPtgxUHi
lsGpubyqqFeRGv10syAJ9dDwNLCYWMwIcDL0JnJYz2dB78ZGnQtQdRgNZGUUo07hA44hYmii6QRS
0+BLGfUSRT3UXhzxef7qThNK78lAfwmBNfrz6fFiJ6eg5i1jOCLfiA9BLx+vwSPhoudgU8F9Km9N
ROrJDOTODeTzgCeiscA97nvzFi5vKt9h4tChGPDYGrpgkg2gDasPizi1JRQ0RWaZ1BgLLddtttUY
GwVn9D7YYWjy/UbfUMifxeZKf6e1q9YYWxARU7Sp34akDTeUBi49t8EmMs4rSbhqrYzD6d93clcu
0ndcAHUKuOjExiFxcb1Ato5+PvnplIaxxI+Y2UpItFjl3e/cyOTCG5al+sH4piZz9jFoMk/l93bP
gNTIAtxabO2u11ReWb0Ole7yCJ2QLbZnSeyxT6/+0GSdQz2WutLWZFDuAuCD7hVrRhJIKr1tom4d
zwONnvhwckXg8KMtpj1kf/oXuBHkuyvW62M+TS5Q22FjRnO84pPuYzAElpc37o80xEALOOx6b+gt
r27o16gT41UxgZDnXIb8VlzkfwGXXp1HeGOFQrFnIC0b1Y9hiuze8KNNTPh+jbQDRcR7Yi0zN0CD
FDcKzZOvpAVY8rlLzRhQ8wmThQpj8vFyNIxsN4lfmyr7EAkHx2uOQVseBc+OdXKI+ySxrNtdC9K/
0nm4L4Yy+C28+q/utcVXYtOGQ1DLA4J3uUzVbo7lhPm4n/PpyT+bPDKwVGm0IT/KNvIUcfD3AJFM
BGUW1n2/nyzPRtSdheARdVHTZqNlN9a6unyCENVwckcAVcd74vZIEGn5ZqO1BD0/Ru/6ZUmQNgmM
2xD+J7mSD3eMBDEYhcRyRN/MOyBXtzaqmcoJlh6FokJ9BHQHLicDB2qHu3PexO1D015X2ZfH1Hwc
ct7ww0xHUs0gbWRW8lt8q+5lvo7O6aUmHM0iE3QLvH25btVRBmrNDV2fYuvcxVqOOZtW8htNLxYG
0uNTvKCqMTa7fGzLwwxmWjiqDvKibRbXy8HEsIAX7C+na+s7kUSewo/Zaq7ROF6kfg9aaoR/H3BK
fl/3UzjSCg3JPFlKx+StALw2kYjTQGVCdyreh3yoinVcbvddXK8ao9RLlZ8F7LJSdu4xb140BFVS
Fg9XIHBuSB/LmyZHdPaaOfnZLXo5UJKJz0w1AF/410W4+DhjoiAmQHRYGBC1x7kqGuhC+FL/EhJw
erqhkwhk8wD5UmethLQJl9LyPfBuzGodaLDyAgmVwYz9C14qdZWZIKM1gQAV7z2XDx/PhhqSuNcf
y2Eo2LYSaH+fc3keoU+nNueXGqVjigN3yB+2s/nmZWX23x8rbW2JHJbFJaYJCUg1i71qA2qinvIA
4xPqcIGE0Yew0Ue+m80pREmao85ehOAPwwYKPJPu1gIz6W1rkKlf3MCmBmQXDtz1fKUpSBhBT6vv
A9XJCs7cbsz19CQgtjxxgxjb7iOSXSsgop1wUVye/eMnlqjx/szKC6A31FA1wFo2G2DPcX95a/Tg
rChus+JCeMsDI+NXNV+Vzz8BfBjBnnnjplO/q+Qjzl65+BYL7vh/Le2I6Ghxx9qG6F1yLTu+NLaA
WfhfYXaKAJ/J9o2UmTKGbdcHORjWJ6FnwkhhSIdMyTzWhNbEnaj5/gzBek5hVgS4GRkQ0qRQyWsu
QrF95qAqkLlLbfZ/OCgFSLxMcQw9WYRKpkKJO3dYgVOHFXE27mhz+tMP2nv+3PzfbutYmqqBTQce
pqWhS+PRHdR1Vs6nMmUuRkigGwMY0bdGpCgp/7gMJTdjMuSbOaOF2v3PK4bW1YjO5M5ffgvGZFzf
btY0pguyYApKnRHRNH2CjXCFRmTrUDrBfGYDSsEFAu7Phm3b4jFZx16aon1saWZiopRISMsNEIwj
EV3avRcP0sKgykyfcPJY9xN/ygwvPL2NVtFWSSG/RZsCu5oa8FdP5DDMHTXsQFEuMj9t0XU8AuAQ
ZsmzX8yUnDbdxx2/+mPqY0ramoF2SY9/gWVIPDjZIQCBC7orj0FLassb80TRQMGofKyYQqKnbkok
6t2NmH58yQCwRei3Ipr2BFb10pNvyQakeqIfrE734YGtb+eUduXG3Dgzv0NxdvGcNmDoo+s9z9jQ
PTCuthHIRVccgUdVJk7ADN+mvroxwz3oKXJHcbgiTLk19A5tvrWA82TToaI7TwgNzXDt4jJYzrHU
2+l7QHM8AC1LM1yRccbvxWyCPGZL2itNbWxD3fkVrHSEiLoTOa0hLXTnnSj7XarA45pdV+sU9Xf4
Zr1QjMCax74oE80tyqfkyCrU3QPYGBKYql0D8XxYYdduxn2TG3wV4yPC+TB9DOhVfcAo87aIDIir
5TNYHclf1ooEAeG214cZu3sOonBKGH+iZSBBL+VH/8PLWt5xn/G2hGeaOxU6zo5y5PawrxHnJrrt
EpVqX3xaJSOXXxpuoYTeRJPGjKzY4R5lDxEmtO1hOuoxHmBB6Ig1OO2qjgWrrxloT+5Uax+1ARVc
w8t9emRlz9lach7X2jUBknr5NuZQmpVb8wMXlzbvUzfegziVncYvUKTdCjExhNG6NXso6dZn/IGW
+CK9uE2lfKpAm7vwKHTLDyGD3qpQhY/7JzwFI96RHpWVPE7Ir7JA2oOoqWNlAGLpmAn+MPCDYEPv
PiJu3aSh8yqYbqsTkBrWkMVwlarRMJLTgD+MKNQoUs2FNf7TmsKHxtJO9oHLh5AguQHKlYWrE54x
0E+TVmFJrVwlw3XhyfSpp4NTzyXVhzXDXDqiH920slWWk2T12DKNpo9oei6LhQMkAdrLTc+qHLQi
zufsH4tu/NoiUeJuHY0/cnDB96OD5F9j/6q+ZBlPQRIe1PHmGxJig9JVUKNNxjlZcJNJRYTDWoa8
H727bO8pU1FH6fSKkNKe8aYiJhPfRblSrJBiqOyJmhw3n4r4/NBoiurv1yFlsI5F5mZeDGWBLYHA
64iNVZ1igL3SfecmdypCjZMDPeNwOHDvi0M5Gk9DhCt8T4VL4BKM6YyODuQjKR5mDBBc5iX4wMhM
5612gu7CBwCBlSEGTyl7ztv7zWMWwfqRHiZNry5dBoWZAexYT5XkUh+m/BGHUYwvd7y2vAkWcZYt
p1UczVUTeoO4IHwuoFPbA/+WKz5Y/E2nUGPpoX7ZCJ0ctyZxts5DwTN/un7VJ8GwqXp2qcicblEQ
hoNnkoLQsSgSM0267kUmJKMUcBiipgEtnn4bX1GPlESgnhwUWe5bIMBO7h1upNybFYp3Sn7cf/C9
Yd0UiIVBhTUPVZI2WtaEPlI6R4bzvHNuKLoBb4yB5czCaJSJa52Mn5y99oS8qGy2ciFa7NU6t7jw
I3OxEpWfHnU+9TlnpoJ8xe8dHL1RZH/jXFrWQO3BlQhg9XzmqbiZKD8jdtK2xb8jiYkSxTK2o9cW
hPf63iDrTnoqxRBuNIaCJDeLmirl2dizNOmS1n9QHdQT+3pK+0Ox3nfQZ4og5VS3p0N2vkVYSsE6
iZLy3QwFqvL4ytz3Jrk19Rax63WEgvuFKfpZ1pMOyY8W/gBx/gk10ChqqNzITaeVKrIUjoK30Yz1
Kd2Kb/WrZtKCWOe25v3hlKJ4QKxAn8V4lF8N8nQJamjWj6T6ZxnynUv2R64W2IMg0gB4sLdFCOa9
OYxJZgIJip2amauY09fiOGH0Bubuncms5MZI9PonhFrwmq4/HYIreLcknHD2xcQ2cjPMgBWtUBEY
+ZmFQKbvIlucxtLfY/g2IhBbdvGW2VkaqbYGHjeIFTG7FnoGM5JHs+9foiKUq6xMpmC7BcdZnrQy
Rj+6lO7wUTa9raZVkTYuZKOTXhAuNTQRZRATPM6y0paIDdp0nNtKuAZ5Yf2wbY6Vn1R+uJxTJU9e
9LJYUZTDgIieR9RH6wMTucvGUFkUNi1m2yYjyTZ5z9HSKBBR0GH9mC1ClRaGmpgsHoXBID+9GFL8
oRX4ZgoJl2tkjhKuuevBgih7LacOFbtbtgLnl81nsZcXvidoBc2zJfr0h//GkPLMb0RUjjrmJKNf
/pQIHVAtt8ZXSICh4olq1q5DlGgzpUEPQ91iBqRuth7tiW2vVB7Jj46HeiWfobm8V7/KP5Fl6UNI
t4EDI+VLXupejs1ydY+BCW8lCAhF8HC4/bhZ45OjIJntIJsqLg1dgiJqFF386wfwLXYBQfQbFDdc
rW0SGAkUooOfD8d/aLuQ20uPh9vaxciLwgtjyoUyQ9dUfVD/LJDWr3lAT7GBZkiahBFdaKXkKYlB
ptv13Vw46p0Sr8zi/83da/OOMMB3WfV6gB3GrOiX+3BVcH08JuvjE02FF7RoXu4VItanA4ejEjKj
LZkQoHF1SBLIlgIUcRxY0f0mynCX7sMgzfvbo1kvS0kTqnuiZMxoxfkyd3s1vPrAIhh3iOIX7d6N
Ly0rYyWlLrhXTkoDBgLfhL8dTWhsTYaNnighHtzL2XFLznjOpq9UwkboHI+vTa9RlR08TmPc0zum
dmUJEStelEVbrqBj/0TG/+E9oGZ8/DR3p6QkJvvdKqKa2/PYjwIo3yIe0Cs4QOy+kMaF+xGHrmgZ
99pM4uuYXcsJxQuyMwZgzLV9Uxu7hFnPZ3u6lqC4M9T815aYhvA6MV5eA32+7BRiQ+3crubDO+DY
HJWSCPMWw/oTCLWsbP49tmGc3MvP1IKTOpCWC+HtwXdcfxeEA+CwN6UEHLiDtU8MsQ3AdeLXF8JN
YCDKHwviU9wM1W/mYokAuQurhOAAYzxZDTgjNjdPgMxirg+d8lLy9xFng6O7D0p6Z9KhCLIuQw6M
mOl49sS5SRC8mZdYTzdZhCJDcSwyFSWeWvSclw3uC/rzULekMRhpIPXuqTjyHKncKLM8tHJ6g27Z
XR/LZNlgYrYeZ8TXdwQS5Mu/TlKieQH0ZUwVHZ6+SWwcmOkFPsKRFdG+4fy/amBntlfHWBBuJD3b
jL5ucAvUqhwgSKK37jC+ScDJ6HUXeT7IkCf8N3UQsaYwo2t9s/Z7e+AAFhZTj5NHTBrUxQFjN3DN
EKp5ep6L3+ObjyicRAMsAIvC3cQsVYu2feiI5niUJ1qrl58WH3ZW/VoeRbV9r3j+ijtY/rJ3CFvl
dP1ppr0YqFzxOZC4yq1JRULOg2Hk6kQDz/35cDUkaml2wJnpbSCYJh4rs1kfjlJ/nwypHlfRCtOH
2uTgZgsZ0ka1tS60PNC0t2eHYtDNZ7qn3BdR6uOtf9R/SZsgr2TsYR9AOeVUGuwZbthdKreRXnxn
2cW3Cs29/3idMl7bic4Udq6ibV+bvAQHVkFYqujlQlMlXfHihg17CHnpSdpk4LBxWhSbGvoJj0uO
CRBjVTKPdOOpcsUa5OK3qpj5nbF4ROaOfh9kuq5R5wTvIsLrXFn76oKmSehcGaPYU3czotc3D30P
gA/ZbJrpnRlrKdsIxC0YNga/r+wB6tYe6LIGfLIVZcWn9mXrOYlLq/3g8u6JRkjBRhcnWy+D3uF1
Yv397FBfivtmLYZldAkD8FX6v7RbPx2F7XgTaXP23O4YozqORXlKo9uYUivrAsJ91hGDcV9fSsn2
q9je19/kADA6TJtrI1FOZBBU9lmqlk50WeiYTvLvtmzqh+NadmjSrfORMrR7oNbvH74p/ZLVTVCn
KfWeDzW6vOMzLTIAc3XQf9q3C0klqURkxV7FItIhBF8YcwVln/NCwJ89VwK8cLABR40tvOWGLNNk
ZQIHAeQug8BqqyIcHh5CCQq+3l+usmSYFAe1Ws2Jk+YYEAspmOyyJgFBJv5XrWtpI+z2PKiyRbrs
dwTQzqp3cpjq1IxfnQ+kqqgeY64FPiUVBVPSuacDtXlsw5a4jXnT5Zf2nD/HORyDfEWC0z+UNBLR
PYzJ1RWuqeXh4rX0NBaDZjKNqr1YTQ9wADIyzislKUeBGZERZLQQ3naOj1o4TRRSegMagh1bSgYm
/CLfuP9GLEQAu1NMTSfIvHp+43R9wrZD2xxh7h2FjCZz5u8/E9qxJaKrvr3Zwm+BaWV8marHzAWS
rYovj24gBCJB30na1Z378Q74/QxZSR9HfCYv+QQowWjN9T3KOhOqg1TdbhLKrfkk6JzKp/WcEAgK
sllJb2BTb1OhUZV3+aZt0566FFRmh9jYPWY5th/OKm08a5sBCzH/MZobQoWtoJjol+Bq8qVHNyVA
dPCtHdoEStRi39UhD8H+hwHNREBjh7Sesvc2/XB8kHA6fq7xwH2uuplCFMIxILV0zR7YKSOMR/dX
wL4hbzhySZvoWAgrJTEjuN4DLYR2s3fwA1IZ86G1H7IN3DI+19J4lB+U/8Jdvt6AVEv4aM0/lSq0
eN2YLPRQc1se0OgRdrzsvNk4ywtYLb+6RlNZjZ6TwIqFoeag+6bia+6rD9kl/bSFxpHXFR2ceyqm
O+Q8wRmH6iB5u5WWmku42QPVFjWNXxudj8SUDVvWA6MslBei60mrBfowh5AQ35V9H+NEzNPb33/G
Y62RNcXiXYGhBq7lCKtoFz/75HHRh0Z9eLe+Njsn4Qx0fyQFOP9HxMJXvZY29BqZ1HB+lNGdSeMp
3lFJtoU6pfEe2swUZi9YjmNUHCdxb8Ynl7JkU3VboGoQtHcN4yy25AzUsUMlubuN/ZSFv6lqlsIy
NOR0C7OkrLny6km6/kqBpUT0bE+nqDRtrbpmxHrSKyQG7SdI9HS3xuGhrGOjlVA4BFrSyGJjexNJ
9hfRXq+0V1qreLUFLAb2iQbR3Cttu6/lGGX2EskSery0ojVrJje2TcvJ47mypg2cwo9cYcmgzwtA
R22UNltEvuDIIrP6oaqFFDQfi7vEHZ1ST5dgSR/sGbEuk25jXlfcYHWJjb77btFAx7ct9M+NJFUW
GqAnNPF8oTDsUkoY3ysrOfe5VdnTVaBhArjr6EPl/6an/ppQ96aBxK2gu0HkcXGygbtXquuC9kbV
Om4029fIf0+VG2RmqC95tvrN0zrzW2W8JDuTlQvpGa6iil4p3H7brH1CD62E+fm7gFbv3zu/iX5Q
BAUoiw1t1xvauAoaMo3h2puXlN+AQXKXpCQVJeslZl3saC/VwyQVC3YcU5byyfSgRjcqJ2uzJiZ9
HD92VNuNxKi//ws652mPDHVQpLLwqd6LaVYCdOk0SVU3z7CimvtpWhi2dtVQwRr9X8Yk+/TmFohD
nnJIsW9S0pX+tVtyU4iw2rbk2JF8ufGitKozEsAU/V8A6hAxQAoIAePdcY7VJkfy5F3gyQtPqRvb
o/gr1fh9FbA4pa+KWOQpvbFHFyf944krJYV688bSGeCiRm0m7ZBLDhD4e8yQZvb0JbnBVtZ1+4BF
lvhAvCaUNeMn0Glotq0W+BQ2/bADbOmmcC546PH5hVKJ/MK7tS24LyvsHA5j9oiJpxrVOXkCpRBO
hiX4/cQmHKkfPFbTACdG7WfsEXtfugW+LPOorWjdnrXzL3RB23NR1t29gw8tOdG9/asD6lI+NuDE
da3plB9mJuLZOwGLJTuJhPpGcOhuo1YXBM2ea7GQE2TiTCqSJKqcyo4WcIWoBHmiy2yEdbSeCaJu
421FEYF1RwSUt54lpgZacy67mq+GLwtHDlXowOItiqHBYqC0y8t16I+y54XAAzeIrTRQnrPMenU8
poCZBGtycLFePG53p18JPWj7BLEYFrfpWbMa2ohukeaZYqPRGkhWPzG60jwK1tsXAJGFC/4zhrtm
nZCOt4H490qfNGVmXzZWAUXBMJXd7a8kZc32G7O8JPDpx8n7EVgnPiAMGzjo19FwZ207zgan248b
xFiIQiE1qXfoRxE1folNqUSN+hqZWnfzjMTelaC2gLN8CFU9/bBQPGfXeDwJcR9q+jdyrE2WNhE8
2uZz9x4ZoiUx+H0t5bjR7cY20x6i/aa7xUdmZpcijLPtwsXMRVFdNJTN8XDFAY8THca7V5qNnt4x
VYHEfrKCNNLnlUBHIkdhZKkxuHgyJXAWA6cUuk6YfuM8diCuJOvSdnnsxbEuyyxSUUDfZMUz85kF
7/bVIbTGkLzwr37I66KA2B3ddnKXAobjjOHjoTmsoQ2P+tH2QcCRqBVtPNDphpBmT9TkBUnZzn0z
i2vFNF9bnvLiG7Nt60khzKPQsylOmgR6suJrM+owVaWKvwY/8q2gRTb+Wj0WeAZHSDhHwNuzFIXz
d0Rj4UMtsolad1ag7lHcbo4q9Y+AOfTa7zuyYPrX22qPrh1KLtO9OUsJoxggUVOzywuE7x7TK0z0
o2QtPzmvz+Ee8pMtq/YXAOnz5WojRFWwvuSuB2JEA/aOeXbv9CUHUDjR7zqDYEsxpm1qdeR8b3L2
IGsN1tjO1Jdq63DSn8GjVg+Cvf7fVj95MxAdcoUfAotHzd/JYaVbLf8TZRa7ZvdUHdjOHrgLHEXs
yd5wyw5j8PLGT1zfvsOPcMd0+h0qL4Mt/spLSYd+exUGvJDfXlWhmOWUepbWZSaHcd8LsHKkW7nZ
3/r4aEnTR2cyxMI5i2CsCw1rxlkiF6yASuFXmpsDCdcdYd9ay7F0E5MUhrDzuU3blmXrbkzdKesf
ZVUGLSjnEqOClVYiaUu55Sx75A1+qbY2FnXMpqDXzpJU6qifdLqzKAO4CUmRtwu13wtSezCYoX0e
2vYfLqlfwl1E6PlwpAO1vfjN1stgrJyqtv/6uF5Gg6n2fb9lw7QkXuyc5hYu4UsCgR1iCVjiqY4s
/Bg23WZk8cb0Jg4+zpnlVM5ZjOCc19ZNB6m6/AYErsxWQ63o6hOCFVsfU0+QNXGc/wBqHUjDquNb
pqk1eKoTWiJB0FnTBu3ed36Ncv1TM5+jg5DGo/t1YGqCxwZGKez/Ip6de6/4blYvat1XBMwmSvaE
+4x8q905LtvCoj2p8/5ZTCHzci1L4Nbw0yZA88ilNWFMrq1G61W8noiP222v/Yy+EBvIkT/ZeGU8
u0UbQhStLmJsZu0rBEJ4S3eA8MRBEd0rW5sXl8J8VtHwtKhpH+w4WV+0YjBeV7xa2labw5xbnTpW
bk7LCtQDgY4v9mhIKQm51NdqiWRlkvIC2XlvhL95Nrg0c/Xn1kGJZuThk/BeW79RuZP1XmL8j5fH
Jz0sFZR1f0lY0WE4JgYDl2cquwJxelNzA8CvJp8Fy+K1KJxgcZ76hxVpGlrolSkx96O4mZMi+Xto
Hg4c0iFTtEMpMgkj3hcRpjkeWOGpr7lW2aAUr5RVYssg2t38Nv0vuljOqsYztLmx77m71kGU0UOT
WqxmNPaMuos7ibhR+c3XleMFYaekTSvFdeLOEmhy43PcOTMTZlvhVre8sNAzFEa77Eqc6zvS/3cM
pkydf4/QNCuF1snU/aQmEKDkrS7AYQErCw21RBpWymmXUV3tTsX5oUEF3EKhZ82bwhZZuG5KWJXl
nosZQZD+uG7Pu5l0xSr5i0KHYCMUYKxhQ5DaFjJyS1BwKfaC8cXtl77SfM8riqtrcr0SJmMGXH9t
gmRgcfsUMdxUsA4U3Oa6BbGl7AigzE7aBWZKnvIkttTlsqtdV/KLjyZp1PqmKDfDKUox1PGnNATK
TwHdPI2EzPPsgUWW+tjhs+E4nOvcrx6UJFhF46XxdRCizLmkrgUxB3GfwqSbW7U/DaGefPFfzBMF
rDaA5zyYzheYGln/L29wUi7XJBwjoGHTUVxkfp03aHcsC8NWm76NzRUjQTqn2VODMwFyMvamb/kA
BI0XhxedH+/y44XGDO6HpNcQZ+L2+iftCyeUfwzr8KJPvSDCmbNNqgOErDXFXK7u1ECirddmMzas
qz9C36fhe4PSV6fOV01z4BViG/mMbCZjmHnLdEbNUPl3+MgjcwbbwdR0pQ+GD3Z66I0tLBylwqEU
hV1quHcF2ZgtBU3Ms6/g4MY0vtaKJMEB4gASsbr+4WwUAorqOocdiL0VB+OMfhHEfBb4ZV9LUyeY
GoFofrur1vMDUj+sKRrUXsK/Wld4BC3pJ/0zG+qTaR79lwNaFR69OXF+6l+EDEmH+7RPC4DvDF96
wTCpEmP/5IuF4xg/9NqnWzKByW1oVKNO2ca2BTwlUQSMWRX8MPGzTEzlIpvQQqWsQZWLnKooq1cx
ilQcYY2vpQR5c3oZUCbY55Osip+6xPSuJqu13/kI36XI/OdKkvJZ5CqHVngRKrnWGwVEXLrioho4
0Z9VkdrFpx/YUr9IjVVWPvPtyfooDh0Bxx+7Ywnb+v/Cl7kQnGnkUibnXcxyITElVPnQUbTwZJgp
eHcH2F/uUSZiqOxVakdi5fdtOnPRRbmTp77HvHBVCjXk7Qx8NmR8Lzps/1wND+imYTFQX5hB+b7f
0H7m4e1RhJLb8AyX0lqFWJy8W6njCa9KAN86rTag5gFLbA1+ZMLCWSgqupORXuqGB5Ewh7f20ZMk
R3ifO7H/951TMa1nVBl+9jTcXUPbkTr4UUjhRFSrku5Azp26BZfEo7IJknfI1+BvPkna4pX0MrZ3
1K5tB9nYEPRvy53GAicUWVrwCpiShVLM15jTLgsEK6zmCPyozuRMUkBd8+9wBCVvFxrd1mbJHhrp
xbQVeqZQQHsilDDvZv27QAbnVukBvzraHm9GDQ1hyaCnE7yBXaFQKsF5edcaD9/PjBU/w4Yh8GxB
YNib+wwFdzWLvTR/c+tY0DpFOYxVwusKOyy3cLyUa+FXOKbwRTgPZ7gdeKgCyEjcxhaWx7HWCG/D
npD9GVn+V5KqS++Co3muYt0beMtx/dR2/cLkBDejHI0oJP4TnIGwBQ7COnqdTpop0/9OXilJx0Ey
M/ABX5GGW2zjdzwsyuAadx7dNoON2Xw84npnatqLDfxmK1oUhvE80i5ecsGAPg5UtIAlIjE1RQ9I
+5k5A50ReBBeKYgMo+5m0ihbm8sm43S5Yj/LnSFXAkhI15VlW9yZo00EZPDfQQuYhEnL9KLc8PSi
2tag+8CB7llw4m33LmbMidNxlM5wUTqvVNEc3xLhEiDP9YYEqmYBHtLrL0jxnbBhT/o0YpQ21fjb
yVCIPCyOb5jiyuagm9NrVls5SIUnq3B8NEgLcrAoGMlNMubc5WcazJqxqWo0z580Rd+p2g2KynPk
utUzqqIP+OB/xTorODwIxc/ttGiammm7BKjcqSWdQtvCln5pAOolOcrZe0u9eA3w7pTEC9KewGHm
opyjX1qItnwneodazH6U1UQekmNIyrlT1IQovqmX1LBgbYSfsfxef4Q0gOMAKQBU9JkaU5tIUQIB
KkcH3pKjk2loO2m3DzFCXGB0YBGqsAUPBsVjX22bgJ73EsRUD2YqAJM2RAMMJm78IQtTYvzYRt4D
aT23jluH0R0U1A+ClOlMIjTFa/x+okg7ZNLzG8hpsV4WCK52QrOG1uhlLx5kOmAF508JDv/aEh2z
RQrrkxzWB9oo6z1fNgJwa9uzAofSI8G4QKd6WciNUAJeauf2khny/4je/r2A0rOIc5VAUJxOF/VK
8RIwE1zMtQaSz7M1gWEaHsYsi8G4T1PsexmcJYNB3T3dv/jy2r5tt6xBywlP3sJChNfULOX8endg
NCw0QHyFn6RT43cf75OmBHNRHo1ID2TQ6pz1NZpcL+ZB41pLn1ti7XK5iHdlm3GJy7Q4+PNhWzzB
YFCr4AwNfHUW17yde+w2AbzhJG99IJuVLC1dvdR43wE6wwTjEajxI3X6uRidfVjwI6/gvajMKeKS
lixy9Hi/sJJbvNolV/Jdcj3b7SgfjtwGvyqhhRpZ/j4eEQpecc3b5jqQGsMtv57hfWNawWFjBkxG
AVsPyPHNPx2jYeFsbM5EvIPVRZiPRf3jfei4EkQA2XJoRnER1UiL0ACpMSu0CDaQxsTpsIJMGEIR
J2RFJWbBJxOkU7TyCDW2OY3QQ4sR/4HrhjwsdD9XzkLbWj0IKVbIhyohm3La2cHmAKPviJg5BTd9
b+DS186t6aFt/4fq9VNnwBhul8aKKI+3jaDIGNCfyofGatXH77mb55bSD1uCKKr6qekBXJCTZjuB
qYaoOg0EC2WI+qLohRwq0d7/QWzBm0upv7EStG9X/5DCUH05vEGdOq0sD+ipQr0OncmmwXqu2FRD
hOFPIVIsqBfFFmM1SiWmqN5owIrAKmEGANsfmOIqhb1ADh72s/h83dcehQ3+GsGLUYcojnql8yGf
P1m/my3+dDt7IfN5RkshO0VI07fouDI7juIfJV59nSWVe0WDV3+YfWMazp9TzIyF5186jmOhUGcW
HUw4UzJyryyhi6Npf/d1E7rqeRZa0+Rcdy1XjckuPVhIRhUNHQOxiAMwqCRl9I/Iu+Axbo3nfWCf
gohUNJXuEUA4XFQHhL55CnsdEWkK1rwOWgrNr1vS5F+dSz+7Wd3nOfjhU+cJTAu59UMIdYw3k99w
x3NYyiTeoTclTqmgHuPBBTCf9XUcwsrQhJ7MMsnJzwDaYeT3dL2yPX2sD2+Pg/O291qbg2uPvo+C
O2kD/GKg/8AVYdVBVNHntKGcnzjmYLQCS87hS4/YU/XYPo79OIDo4CBVvtscZavboGH4H38/ECRa
GC/xAIITI6OT4j3ugc4SObRAi/nWyrEQeX/LEe0HY3IwD4sO5TzRA2c8O4S0zdcSTW/AYhFdYC8D
Pu46AGDsvfOGvZgcaGNkXIQKqQtQ68fcWFZ0o/HmE3QMxS1WLW66+p20+tIbfJEcQVQYzXde5etQ
+tr2RhKdeboLtgLPQTopHBvzNOj5Sfl9QwePyERJ/Rd8gzWcJdR+QCumLQoep8UyFt+Jpa7YrJaQ
rQGMsBRgVCdT9ZYYrTX3HgVb35ApmQJvRrVSJGchQoei/j0L/PaalnC+2cNr1hWrlWkFO00+faUV
/ricLVbfW+HvAOVifJzbB+KF08UI+VdqeIVcp7p29PUSTZrEPuFnTRLkZfvhKeP4PKhH/Dykzy+i
BHxjaa5B7Z7pKkeW9asNqJ8GUS3PdbIE7a28lVriisLoVsKTQRDUv0ud6JuhhoeqRku1fMGGkRKR
zNkvlMkqORR4oKt4ErgIfLSJFKtKRSPwvul49kZynQh9Is24kv1mVIHzTjlPHi9v3H3TH4J6vSpV
M7dHrUvXLGdQ9KI9k36A09Qmuv7xkeTzNwlfjyVTs7FEBBHz2KOeEsu+ydSDKsT1/yAahaENEDiU
CZB7dErWjWArP2MJbOqvFLe9gqz0/A2riu49gxUzH+A8+UK1xRnMrPHsdnxswwWcRGnHXeDVUl+L
BUrVAaajpgepqUT2bqApRMWk7X3iO4RgTpX/lvU5b5GtwP/jddtE5203vveiggR3L5gw72QbY6qa
RCsKRb273TFakhCBmDM8FuJCgOdG8ky8CBIqiduwC3w+HjSbLYnWgHT6+/mERVAxEZYu8dk6ovFa
cJfXry3VQVZKqlzT2bl5X77wlFvpdvFP5ADM5ljrtH36+ib/mA2FsJYwXQAWcrV+Kjc4GppMA4mk
O8c3uGUdgTOxInOQhdF54I0IonlWs1EHbZZlAnJP6mrLFn/8udWr2Zi0kPvRQT9GF/0pXx7QZO13
3jyuznP8Z2jrzOfQ7BU/n5TpGaiQpyB39H9M9RbuNHJbFjuR7OPAbicuSracehB4mBeZQV5Q2VJb
+UJssEM/qfp+/WQOE1dRr01VaORSaTtnIQ5psKLKu4jOXr0fLEZN/tLvX/Iousi/y5XsE78h9RrJ
W9qqEIZ83sUfZB8V8Z349NX5cUnGN0qulFIxw+LFnXShLLTyeSC57LNwxtt4sGk0Qt+icIxjsMmq
SPRcrpacKj8qP3M/PRQrGLUOroPTSpdHb/ELE87X8qlzeBtnzU+C4forgJptAo6MA+QtfMR6c5Ol
3+sCQSfwnkk5y9/LHvjs6rpLp4ZV9wkrOvn6MxER4KJ2m+df8ixBKwqgydLBQ4GMQQ5u+s7u9rks
OpAtnxGYysDgl4CI6kLjukK0k9ffKjJ2a6+SFgyHmfqEeXzqNllN43SxM7TnDMf+EGXKfQlpuRco
cyZIq/2ICf3Na2J/zkZjEIrfbeRIVrW1HXx+uoC7c1qlbx4KgSycv62ESd0smmdvW0/4/GFn0w99
/hjTyxvNPQt21dtdq9vjMcmTWK/z3V5aqlLOf84ntBTK+ZVtHkUh1nkuzUX2xiQAEx5mdXbmX3xe
/sQzx6AS2FfD9G/rJk/pPhkfJh+I3YE7KAZBLbG/svCrRqM+/BjaIx4xfZ2LLbcjF6cv69Eh06fG
rV/WXpMTsP0UpgkA7ZB942NOETIgLMVX5SAZD25HKQ1lE0wtV8MgM8qUJk0tRdurk8Skxw1RtPSQ
BXmffQhBYuGLneeRpFjEadUyrHE3DzivPT0csLg9wkimOns0Cf4hecEaxsBGAAMf8MFts4kUpNZv
UB2lcJJ7d0y/aSxia/1UrP8wegmyzanBFvC9QVz/euHTmUtVjW3b3S6OSiux9V3LPI0NwVlvd+B4
5Gs8mxcfCr3bHEr4Imo404k2oBv7Dzzu9GnQdqsbI1ZgYAMoGRYtjvXuww/qI7peNcBON4RP1Llt
Bo6iOV6nbBLR5CzSuXRDeR83AUqlfBElgqzPwUmr8upOcDkouwGadsJfLGtE+XTgbswoY4UOSdfe
MKy0xsEcd2GD2bK/Z2pU5FDGin7h2OkV80N7jYhnurGKZVlJUnUA69f8azQK97uQANU6rIF9PaOP
4ijHYXOwQElBZOAP0WSsSeB2NRQMYzvZ/jh1igpK1AaiyCdLTGyhJAc8eJWkijFs8c540MUvKAw2
99Ttn+wMZ9NvVTpBP0C2ADX0I3tGupfhuLroLAJ4w5Hp+fRA/5eE2G0xXrqmWfML7Zje83+cZacC
0WhVosGgiWHz4mWhNt5b1WZa9inSvXJVxreKMk5IpQ1ocpmGsEgPAXSv3AKIYdP254CuaBFLCklY
lw7KBHcPleXBq4CBlsbd71erlQtnZ5WGX56oMBtCW3DwSuYiLBiQe6Xf4JFMXpYW0de7L+z1JND2
UQ51lab93DD16md8LQFXnIABR/9P9xwFcmZNEaSzzYJMZZWA77y8eVm8DAl5TgGZlwtGCcW3XggE
k2oSLfx2v+w3swyRhyhXFLIzms05DLlZCcY2DeAVhbNrdQgk7l4MBX/qS5NXbyqX2wpmO1FEfbI7
emASopfBPgRnPA2uAbM1ru3aNZ+U99YUS2hXCrEajpdq69IvwucZU0XA0WPZVSsvopHLjdwYkL5U
ZergQWO3+vImxE0HUyy0CTHOLU86DZkWSLG4Z4d6wiHoXEiSqlmYpX2sTqlOhcrkWYvwa07cTTKi
foadTaESx+mhqy0WbaYi+Odjw8jxtd4o3iJHCnvmgMplVTAkT4ebMbC6U9MpT0MMxwIBdyHLt1kk
boBAiNLH1zAkOP1Aq6yLJVWGTFfMnyryNB1lxCYZcK3IcbUOahOfR+XxB6sYoQ7EvujKBN2vkGPc
VQABifpj2bnD3SPLKZCSoVMRHssv+550OetLHuj6tlWU5h2hWaU6Ef23kBuxn5h4L+ycwcaC4VJn
b18s85RFhRlSY69Ah1GxYS1MtRxevTTxzoB/A7FRk7xsePllb5EXceqP5YPZ74KJw6jSG1MmbQko
XyGxzJK2N1atvp0EtDYzvkqIV0+qHme+Ydajpkq3mQWzg+Eh+C1GcSUxFUXXb5onpKlrP/7xwCFB
1HgJl8vcfP493sRA5kOGAWibqJCFibK8/8qPtI/b0g06d9A4SXOnv9VZ5b47hEnDbcFsLLKcld7o
jTvZ3ylGdKFifQ/IVtvcpbwXGxxd7BaciTeQvzvPRfqjA8pzEDXgxrTeaGXYXqzN9HfdlYLMhGDM
XVLDZ5nN2wBCq0MeyJhLMDGEqHb0bXhlg4bjxHiC2YzNB6CSZXOcglvPsoND6vPQAchuiyk941QY
vRldeFPvkKrQsahIxyq0V7ZHAGrXQiQfnSJHPyvtA0tRSywuq2NIRAVVesmu0vJm0oQ8fRLlhSAY
GbWFHCO+4jpdJc+BqJ8we46SCEoWNCmGBnp2jel3WzxU4mjzNAVQKDvI0qQdQC7rk9QGABnZsmys
chW/LQpjPscgLkuAlKEoJlpCLajfxbYrgZyA/QTeItEIqRnVIlju+Ag1ZkhGAjW+4/UgwrZ31VcT
PQ/xrO1mqM6No5zknhEM/Llg7Ye+v6iz35/m2XdAf1QPF/WK1Z0VE0kbdBARdSYSm//o9f96skCj
r7WNLvHxsm5Ma8AJdNuU/fCuI8deGPSRSx72q+dmhWSMuvvAN4zimikMjLJGaagEEdmSeMxRnDIa
NZEql2l2uhonVHV1GKO244YN0y1qCPR7ZjECtdar6z8kv261gXcgdccbeRk0rCnn8lIOeD92kCSL
Btbf+VnolWZbfv1gNhk02AAx1yXtq3JOxuuZs6kKj/VYMVvwuXpbcdgz2/Oqel4fXOgAjDmW1+wM
vP8jIit4Zorz02p3Hr2n4t5+iIrWvzHbbABv+UUBCyhYpxncLjLJFnBiSb9l6WF4DHnAmwOLEpzO
4b0JsoKZKS5bYr0XqQQtDPfJcgjw/peyzl0WwEVKoFw85osugZ5Mszuigsw0HuU2gB1Rk7O6JiJT
3G6APStAyPnID+fUY7xxuSvUabzM7hYUZdSFXaglBxCgCRgpzRgMrWRKLPmKsRSmWgni3zdd2t9c
63Ur954IyqtflBMJUegcJ2xRdacXQcAeg1ApTFNJE6b+CwT/ALHQFF5mIMhAPLTFamN9icb6z5KQ
Vaaeb6YE1DAHLITZZJRimOYqyAJDTyQDNs4oeRaK3HzO23B8VszHNb1sXxHuy3jPosWxupsoQH+k
jlngVeBmkd1B7X/H3NBDShJ8jC8WfhGPMxgxl8q6tOPNSntr2tomMV9/p0AFXV+f4i+Wh43Y00Da
ZQWUkWCSBOErGP11knHCm7WFqMWJYonlGISI+K48gUwinWEI8GwNMncIa4pMwYDCHcj/s1xmsYDV
7XfIkVsvdqxdEGCq3fb7SfK3Vdc2eFAiQ/wK+l4YZYkr/OL7GP01BlpVxmsxPf2dqJWQnBKcJOaX
boMjGNkREgejxI8HA7Nq6tERCml5/5Y5vhei6XUudWH3aTGdjou3QhIKhTtrs2K9hohHgcUjCpGZ
FfbcaoEheHJLehiQ51oqsM8CkcpcjUvajOufgG2Nji4j0a54qDzlf34Up8/X4IkIi54Iw855pRk3
0E7Y0w180Lr3ZXBaRfOmH+vWAw0g3vc9mM5sjSIcESKIrURPGATuc1HIGmPvCMKwG92bdrvJBj82
aqJksMWYovASXhwqMBnmOqiVNb+d+XUfL4Kg42d8s1zwHWw6aguS4prXeMvjl9lgUpG4vten7G8m
TOyketcwaBPvG8NmdjvRUOOlvHcOzUXcKltM0nhswND0s70KEdxQQOsn+RPOlKqsEHRzpTO6XM/0
n/NRoO0tprO+2XjeYaYeWIDGDh6BngRQ13kcCi1W8WZQbIUnKvFQtL/FpmQo4dnEWLxpfuMOUXiT
AGC/kPb8R92pqJUSCkcrC92K1Vo0WV3xvbFUv5x2UsVs/8w07/HG39+mqVzPhVJABEms+5osm71r
ihsGsDqWHEJ4LPWZp/K43pzxYYmRtgCxCcMOAoLR54xLWBo0v0vTDWvtszu4lVtAU/WQj6m8GWOH
cOmJ6a2OSsuKxubpPrZeHxGVAOeuHLyBELAxqbFsU+l1/c0Ap2VhVGHxUg/HJJsXGEZ+S2c0/XUy
feerrwfU8MSSCS5WVR77A2Or3itr2lSex09+2MTK1GjL0r7HHkoyVUzrSCD4pL9mrN0pENOYE0MN
vX1HLltCE/JHPFN/B9C7SD2pzP7QE4qUNBOurcdkBvzmjfPvKZqX+hwoGwSQmunCWT9A5A9izx8Y
r+ljhb8OF4NN7XmelQUKsNr1rJOJ4QJqg3+uJDd4riRYCUcJVtQdZ/olIAVn2/z0qoU36p0CAkhN
Aap0H3srFR/pJN3aytpHmxyhWCd6vDrV3CdHQ7L7p/YiUTOT7HWcf4NsMUI5IjZI0meEq528FYXd
X9iiCgsrlnwM/+8HN/3n8FZRvRK26nus0hNmQvM1ojtr5LyW1LDt6zmRF12gvwMSVtV18Pym9iic
aqkmBZzYaxohPxbLrONbToezmutcfzwvRLf+coJ0+9lf+7pG7A8lL8snn9SXjvb3qEAgX+1xLsKH
cpZX82BkbwKhitOFcH076GRxU70GmqfYy2j9xATui73gR0VsvynPVSosf2lbNGn0PFQ0MzcRr82a
ZJUnUm4JigQhoOGqYjXy6Hxh3BZiO/a2V0tsjgK9LwY9SBZXalljEKZrNM1oebSE8IK2kfokmglz
aILDMLpYf8aQj8jDi2bpZJ3l96MmHAymP+zY0//FpSVhCGCBh1rKFVHmlukfpiEUWwdG9gmyi6lp
oq40q7wOeOWMKlVeQm2w7Lsw9fYhMlr5juRz87OeZeE0EhoX2cZQ6d0oC6TRqtSdOGI3kKsuzDB7
GMY2O9b9PUKPZpigHeoXzXhOBJahUBG988pMoTYfahDxcZ6r7f6j7md0VokHSNTElNzQTd13Tb59
Qr/N3jNDvXzqjrNjDgFcSIU+jIuvtY+33bfs6nSMeiNPePH9iG0Sh2qw+hapd0Q9ksLGRIT8fGX9
oXvssxNJWvOQaKq5mqIzXn3xibbr8T/giBBs9ocAwgrxO8CcMTYiLxPKTcsk6rerAJi9jmYsyNA9
B+hfqI8ap08vIZIeU14D+rSrn0dE18XAj7UngML9nSm6hALgQePhm9lj8mcofuVtvAL7rTtUEq1e
f4RXEBPtKHQ6DhxAe91ZlRA7ru2QK4Ypbd6xZVEl5ljWCXEo9gbl24VUo6hHll/n4X/HCev/dWSl
CJQHwJZHQwail8VFv4pBHwQJX4TiiU2pR4gSmnZgDRqDMs6a9xbEmL+ejLzlhxrX5EfyvOLXSQzb
tzD3hdu0FwJMM5YvsxGp8h7qS/JKkjp6E3I4+uu/HyWbHGHZNBiX0tHhplgtTd6F9MOqXYfUfdhj
5tCjGUHny3R3h3pUHpFGMem5nZbFs1g6k2pGFOfIiYcFuQfpASahnMnnrYVoJIY3NfJbcPhFjZmq
+2qJHGwQ0Ld5ca5wV88FTCCY3ybhhNfpa4nhFK36ri5ZEwR/AZ1CVv6lDOPOwLL824UqMAOhe/CH
nuXlCncD8v3PHYU3YU1pLUszLQmfi6fdeBMoA9R8BfaeJOQ2dIsbozuhbXW5y+YzdHxgS3Znm1RO
BsmzwukW4OSO1TR28RwCIbueuWEgTQ275GyV4YQKplbjCQGB5ICAfPF0IB4CeqJxMFWQ5GGXbDs0
OProjU7cXP/LvZ1dNOk0E1jpbYV7Q8KDaND0hllLBIEwSPlxLwUevydOuDP04gZieJc3UnBO6gPn
eJOOZvCyDm2ut1RTpPi2Cre9n2oHt9kjO3ENPdvf3ArWkdK6yd7RiePrEMI2OXqbzaNT8vCDLDUy
6X8BBEzdASO6JgwOem9ayMOvcjyPBawln5/EzRnbiLeItT1+ioUQQlzwaFPKSC326sokCyex02Yi
RilLPc/p/DGj7iZ63Rfx0o3JbwTQDJaxdxJfNomisPLHwSITEj9foR4N9ywmJJ2jSlf0GQ8Fphuu
EoxWCXnuJpA4mLKFb6jkVK3sNtmMpfTjGrhgOB6ITehhFv37/UbP6VTtla/J9iF+hu4zo1lu0aSS
4OJGf94Y93ke00JzKid7sPFK17JS/FDmKZWjGG0NZh3Rgg4dVOZAtE9DuRClih6L9WdjVMvLfCcH
kcNYObKeY7DUbWNmTVVqTibeFrFZwfqWsP+VuYcznu7TGqM7Gwx5BjpOGHI7Tc/5HrZQ13Rn4SbR
7UUemy/gUp2LkyXAo4E48NALtx0eG4ls0X+8k97TekyqweW+UY7upDxKw5RLDPUy0fFAaIN+f10w
ijYq2uzsRK2erwHUX2OY2mghoKtwpqEZuZpgt6auh+aeko/c5hIlX4+VbYcakIBf5J+eIzc2gcrj
gKzPdqjbyt2CaRDxyBaggcZ7bbLC9fVOgyghHfVwfxa/jt3Y+SR677MJfx1FSG0rtCgvQIpDaolk
Xttl6UlkKqxXj5GLZxceN9gVBaHbE2pX2OJ7XPDO5+XTWxjBLE/h0FR++E0lSGDmNcrbVkM5i0Sh
Z42zELgIfvzwB1qhcSaApDd/Eofac+eTF5kbGzOdsaSYbYpQff+fyd+hTkxHV2BlFJzN9yKScfBh
tL49o+zKT0VwHfljemR8wwqwcY+l2nAyaFiCCoKkqiQmU1bWR8HueW13QljjjjpGSE+x1T5DzAQw
WgFGiGkaMl/aWTu4I7mRrASPY7vMG4t2qS/hSwfC2K2zBuSM9Es/yhocAk7m+MqXgOBW7OanfqGq
nf6LGjvmAJoMoLFABdBRqzH+w1ym60gDEq2kYTO35KGbWhM+PafHobgjLGIHzaqhDEh10jAOutt2
R1Iexd7+TVe8q/dgvFsSaomUYGj+IV5sA0NKqZsqpNLVvNej2e40yZKrZHA10PIMDdRlf3nHUJTW
vOJGANoFlEHSZ/GWZtw7pOEHcp86BO4sL7XAlnKBDp8GgPMiI7V6V8uqUobRq5lWJ8mGQAFIKqZ+
/7kBZJJ9IeY5uLs445JsIVwv6+ml0IxwZ5fU4dtXOv0of1X4pQxruagwLTxMB1EX1qcfB4WN+eg0
ug8Q6qVgklWS+22ab0/JnWxt0qYANwqUFFrzJEy3hT7lLyLI0DNl3f5j8eQWq/mBRUwv7IJt6b0w
zfJaiCxlXK9tTe7YGXrv6+zQwdWoi7ZDD2pXNYoE+GqIlF4VdZkYIgWihkwh2eOpRgQ8vhUD07wK
97wxVq367kafuPRxZ3iQExEmCXyTsUwcyOjuiNLprQIF9x8MRIOcYZlGdALbp/DPFpxB/2dOFDPf
is1r/jH0IjcEv6CdoXz1wAVBfuu/qBM2tqDUWbfcDDsOavau9YFpMhLefGtyMyo7ErCjHL6Upk3y
6zNey3RaYmbxJwigKESZNNQUNCUxnhPiTybBDN6YzQmF4gAwOJcAVwsR/JRdwfaBZ/BiQFjNWV/c
4CKMcixE4tPlLk2JOieAVC3Pbynr8JFuqN9fB59p89v7he6yPAdoj8JNk80M7U5oyXO+RFVs74Qt
twxCHmBqZdQTyaoTDGLSJ+Ur7dbi76cyKFOlEABEIelVcoXbdRHZP+zyUDdnEsTpui974m3wbdK3
m2XeHJL7Hb17uY9YKitG1Am0cAfElCWRBOfyIMn9QryMAENZczaxUS1s1o3k5VAmzeYBtzdpdN42
jWscmXqDS7fo9wrg59Gw8doi2nzAro3JnnG3xEZfRk4vMrNydHEsJb5/IVko6yS3UNmrLaf5Bqlp
+6ftse5hnRMT8VQpshUUWM4lc1Ah8qlz3d59KtbkkI90opYNtFK+yp9irXYS2kcy3qwAhKq/v8Qc
vJ3ydHtvPBOaoIznX7kF36DYsn18b1J7epGARey5qa8UMEaV93Am4YcXtTBmJgZYLaVxxUkXzHz3
SuDPB6EUGoXG8HD+O8abO+SWrTE1kOoMBbXRE/nDptNwdMyEbUDH5d1qLbPeZBNp5vNi+fKozCjx
6M4GDEQ8LwJq5w1v7DPCHAWd0mtJke9y+rbYAHn7yTV4TYw9HUViMx5dRhhXxaYFBOriSoBi7dN1
rz0KRmDj2kgjumUz742R9ef6cDiqbQiKUJ6kGMrGTkZEkUfhKHbf6V8liwKlS9cvGPHOLqg/CWYU
XmsxgtLx4qH2X6x+gzTPGLWjl7XaEXTi5YRkqvcpQKz9kwu3CEePFVhIYZRofXsqynBRUq36D2PA
L4wNyZmNb7+36oSByuiNB9+LsIOV0pcghsle1pI8gxgpMGVLdoTuejSgHAjowo4RP4YObgwYwYWc
4TMCLrPgOrb4kKPcSZ/kiLbvtf93XwX5ZCMAcoMyCs4tQNjKe2lAxyq9n53jwLDBS073jwwuvrM8
KEM9tnucIMzpQS+Z3m3fzmyq0LZMqZM5DYCtKQVv2TCWkxXZbqADLWZiO8lE6KHKu4EvlgbzVrFH
KWuSNKKmgcAr3qa384tckVvGkLJ+DQvdeuDbAfGFzIZig8nHjZOV0Sa5/YCO2fCipQJWYJqxi6Bi
ZVH35z0dBgnwY6oDrFVlPzmIHhN978n4prKGrF6eq8GQ8ebgFHGmjcCbysx/BrC4Bwo+JkAp3yJ6
gqiwLaa5Y/MAv0gvIWVCixW2cNbBEzYHYlu/q2HYsXLuNc16GLwg1NtiDUPiikAGc9zxIP01JvV5
HX9a9VX+bYJbrjW7BX/NzGTk2N9oQPp1vm6/7gEAyCo1CwggDcQ1tgOPC5b+kiZEkZoo1cSzmW4G
PV8woQTo+Uc6KYzDxEgp9FxwigIgS0N9OteQwtTOqi6vCzTss1ZRHZjeAiv0fyanJ/bxqgQPEQEe
7/7LS2xFPNkF5r8Ex7tSG+2AXBpPwVGr2bb8IHh5aKUKx3hkVdyJ8l4TKfbbroVfJbSGNhWFETmZ
F0mVNjlSlRLsEV9ZroTXbBD20eMTQeHQRjNDlKQw+7fZ2AVuIGJ5/jzH6Zf5vpDF02BDKMlmn6jV
KQfOet82a2XTsj8YTt3RJgkF6i381+sXa1mjtx4OG/o7RmJBORZCgYw16fTFK92BpudsEhkQmFtn
q7friWVxQcp+cqQOBUZMUBBFcaS2vl5BVEeUkOGY1iGCy192SjFjVflhvlmy+iapWODCiywTEKb4
RmE7ny9V8JVZKQsOPup6fCHdepd00neF8DNTSu651FkS53zJgyNlGsZTFQsjX76e0Vz/hQ4lCldM
qBZQI+jR5hBdX1NQ2jox/1zxGO7OnMJq8KjB6vu+7RXPdTMYL/uIEYUudHKrjqid/j8WIETpgKd6
r60pfyi+WoyR3Xf1sOWK/AQRWWLtPr4Utj2gZyuF/oZLd0F6xocLUHLZX+R0knzLr0tpjwFpImTc
fD0aE6JMEBKGxcjxReXUw9fMwGaW77gZa7Xbw79OVMQzIfJ5v6xPnr4DNVrmTpdt0Vy6NkQZsAuG
xBMgzXZpnn0CdkkygH8q7cyZkmAt1/mbwLL2DWR2Xq5pDIiC5jrunlSg0GkyP3t1oC/3Udj/TNxr
e0lhnFc/jvSODTCyfgvmzugQdPj1RtN/vNKWwHdGjVuX98x50t8SIqETLZkp02pHs14swohebrPC
ttze8pY++d/PNr7ekxmLXPJdmXbHFaFKJZQJ33bO67GEfv3CXaKtHmeXxSl0PRK2iLDsmfSOouv/
P2tYehIY/cwxVqKpR7Nc3fPwmgvJxLgsrQz2ewpgbu84CeHxT/jBA83tJgFjYxtWltgFCSRgrhUW
aYSitQXZBRaTvcFK8ejJ8vkdkT10TbXb4lt5TPauluFWaSm2y4EeKT0USmbrtkf6WgFapcqwMJ+3
RzpqZoG/69kJPMSFriNDbCBq/kElKRTkcWvn5mPm1Xi5EQUFl0yIiphcmehWrTq+GRxrEsOtWyof
IHJ7VxQlUKOygqmNemx+nj3La/7wjT3ESO98yxH2ErDO2+O2u5NVgQkKZNnHHdTsJijsbAoccmRK
xY+HjbtP40jhCtuh+tz76tCshjf309jYq1NFaJRN7hjRWLG3szxd7oT731LkhzOgl5Hhv1SKkz2r
N7pSU9D78kXXGWK2sRZeSN0L2cPDxNrOBDVrhYsyrYaEkmzDhQE8UxR8G84pA/yKOH0pPPSw48tC
9qn3vFtm3a7z1Uy/kXRQ2MFD/Qj5P71GR51yaLhu+LlhwpHmm5rspJzYuWe3dSo+aylRyTvqD0Xn
Y0VHVLZP0v1i6HyTDlo5C2+3PVDQc+juEuc0ZSbOYF6mtMZpv37BXjqoV5F1uxYIyve8OM3CKhXx
Uo/BdZB1W/vnNacczUM+BJs7UvyhVSsUdc22EN+l2wKyYtHA3pxLlwZ0eUPo+VfPrdA2xJkxhw9/
WnrjdlbA6vZTuRVu/aZUcga8bsU7+otdp4J/i/jwfmREgoAhb2j65VJp18YyEgOlRRrgSLnR3LpW
jHQsmtgedzQj8MVq7kekb4eUjKdbvoxy+KLnpShPU9Zv53AQ8dfT6blozNsyM56BwZMWO7RjMexJ
cJ3Vc3n38iIyXnHRva7ZhLm6grli3vhs/5rJIWtQTVpssH/DaCqOy8C1PX7D0QzZdfFg8Mmcj5Bs
xwa1E25Z7A1F4+vPYLGWCJ+Ho4eOtEcPB0TpmO/X6LE3ULFEfdunykPASO4lCl7Z7u4bB0bkR3sk
yf3kX2nQnie6nBOyPXqOiJ2ufIxxL+AFHj8SCgMX2DTpzS3ofTAnbrdb5VhGxZ+QtGAo0RWZ1L3W
dVzw/uYmpCHkguG5N//CIGeJOwA3yoXbAyASUWyyUZwu7wDL/vAyzrkpgHrKQTQjY/dCa6iSrBZP
P/1LqJ2sKSqsjy2M+9Mq/GezzClih0t0wO3S53/8+se5TZ2uZVf6b3NCis/0bPjDldDfhFl0gls4
hEyUVLTOCEYtXHFUDHwKYzXRfWU3hQ5T7/EupW4F7Zwz2eu3o3khprRLnqN1glHzVNWa/yZ1Nadm
Ks5sLNnD3Bewg/tA4hJ/oXl0pwbDGWP5YiFZZ1c076MagpkccLqArU5Vc9tDYFHBZJOIhlQQgAC8
M+4a7t8pbKGtUuIw2Wq/u/+T6flCFV7NJwVe/aSIw7I7os8GxJURmDOcK9Rp80bgkuVnH2VOpEWz
lj7NKT7+JmC8KRgJFoVpmulaDZNa0KpwJD3tEIb72Dx3GsxevBUi34vi8axEqE7SIMndk47bO214
HmMRscz+w09Li/8iEBSv5f/4XnfACjgGEud1kjSG0blOsxRdjd2mDrqhJmFH4HNLcowgTsDm2Yx4
MNUBprfcapaWQeyjFxqehujBftFeD0pnQYQevk46m/DDWMNhXENI5Dfqz7uK8y9HKNDSSrNKDWw/
APB+zlvIAcdMZ3Fdvnh+Hb/8iRcosbV1aALh1B/z0/BnfJr3vRblvixfJsJlVksnSaZSsk778KU+
QVJIYMm8hVPmLM3vzB6gKh7pNuZNBxLmUsFuNEDG3skuIFJwS4mwWTofmKeJAvQCxUJ77oVcSl0T
Gy+kZvCXSgzelowaZxYxwnmkgFAabTY/7X1UnbJAJZH+y3EeNXIDk9AkV51nN7hZbYHYGIIAh2Vn
hObiRHKb4B3Lf4Pfbnfz01wC+GgIT+bU0DTJFYHO+iTK6eaxtybY2U4XgffagbdL/Xu50dPvMqD8
MB8AXFgmX5cl0R4j8ZYWOBRKzloFaxv4xOfqb4XCfDHPYTek9lPW0gk5ao5uU0aRr2JhXm7RzlF4
HqwbW8s0QZEMM5cvySOs6fsBSQ4SV5kAda7btGkY9t5MSjuq+k+jfex3J8B3Vwd42ZanpwLFuYVP
JIx1DTxyFsGyUyY7rSQ8BYjH5FID18upFFyXkbOeRYfW38vRsLI61xmSJ0DjEWVnI4fBZLMZ/3mL
f4JgPl3CvZ3nHAsviZum+h9QQALNJ8nt5Rx2DEoJOFtcsAb543fv2YKNLlp7yGKjxuaJLmEnkTGc
oLmEIGJcXEQy3Qny9SZJ26DKEJUoS9AqysIu+66LWE4pv3JFuwV6am9Qg48p0Y8WatDf7oQqrstq
e5HvQTWwcZRaritMRbB42dHDQuHnpAGjTZ7oL8wqy8x1vcjwRkGS09w9MHnkZcW6cG7AQGiaUD4I
CgHLNcHtUYTefZfrDNMGzdsn2efiA0hxgnj8KHOfJfyvNLkB1McfDHrGtzKQj++oc5Csb3D7uRb0
8ND7b8VWd8d7K85DJSzjXdUx3Jx2ztTlmEQc1JN+f7gcGpd6w3rhNmVI4UlxeBozeAwE8si9KBjI
uiT7pENDyibXtpM98vj0+65uDlpcTU6BMGvw69oPVswbtn3vRbTYSsI3X/PZ3rGdUHJXGAgNKpm/
idmJhSFglTkEsMZF2PNo+QqgcNf7LbqEheEfPhNf21AhSMpA9mleKpvaEcxrHOZVXoueU7hOvU7h
73gQbSH2OKsod/n+fNLQhCV+HUnjmqnr9v4yGfry4tXsODbhOUTCVzhAnFCTcLWUBQXSkXVejH6O
KkeBmE16mUhxM6p6clkRyMbZu0/7QefJ8yc63SGI+d77VwQcXfitWXkRZRxTJzCyD4DRNVdghlpY
Pio3Y+Pa2/rtRNu/WLocw8u0V37UmrPGqHO8bBgKe0C3ZWFqrmZxTy+0b4lHXVlJ2pBCdzaaZTJT
IsumpDGjmEYs6C6EsyGYTsLV+JTz0ttu7A+HcqOqvhSaCBErlWcCM3BJ2Upc/KLi/clQfp5rjbPM
0JBgNySHqNDYdHa4nvxnUrXPqIGHT1REUeGYrFZbTXtV0HCV8ndkhMYno+s1TJ+wRmr1y1AasXh+
8WsvtnY2sBsck2bt07wJDbqtuJavD4ShhpEWnzBVoauvfA0APMPTUw9UrhIztpk/hdrqJeNWD9g3
kr190Pt2PTiibgz5et13uSt0bnzrSIEk6uyxUhvcx1Fxm4wU5jS5cq+OIycKQxwDCFTHfpIhlGcO
PrmCZ0yRsVMkUmKL7UZ8ALE6HFsJCxelVsu/g+IFgZrqT2d31ho1cV5c5KlihhwznPVG6JeJCY3G
/cSkVI52AuPugsfgonvbTGy0CsJlPhtDucfvB7ysYDGko6g8VLbA0NmU1LOxNXp2nG/F0DYxoUIR
qfV7UtMc2EvuGSAvgWXs+lUN6iDJRWXo6H+3KTu02rqODIixtrHv5a3HjEcdORlLoUAsTnqDIXHn
FDcOL1jQZksIXuNGQtWt4QTN1WrBjYGfRij3OfijEUrL6+LSz7bsPQRZEbiGzRbKg1XAy20YwuhG
gws4FhRps7jYeimx9xsKbh4kLkglNZ7yxa8I7LunD0P5CmYlKQWiU1UbYi48OtKxmFwVo+05qJNo
FeXeLmU/3F6NDlrv90Hk7oJHEhKFZLAySG5HL7W4PgRyL3/I2rD6hgeOfmzvvQJDVlqbM39mDDQT
pipV6lepJBkCTFawkSdLr6sQtplsw8dGdhPE09VNXNgORXU615NWEgQl9JARrSQjuLx7InmwcwYJ
3Hm6rXKgSQsirLnbgixHZlFrptEnIa6G361uZ98H3dc+fWclFkbZGYj/TC5wIBAnBp/iQPnUuNGW
tPFEutpam0S59PwmUR2LLfHzG/FPuApkQK9fvy2lV8vOKalueyNCgApvEkf6lc0qSw1ZYdEXPkoj
KHpbGO9HMghJBJgtf65xXL8l/IyoLbTVfhAfRp4trRL2JKGbw860cexQBLoKprBjJ64+0MEu25Gt
UlTP8/XWHKXVDC3jEHHJiqEVbhhdPDopo5GSAaYCLQiskU5qbO6digWopCcoh5zQdL9+2HkQnwuz
Jp9Oq7W8QEOM2s8hB6sB3edzz9uXkpizJGmY56lyn4HojoUM2PjzZH5JnRwTlGr4tDupfOb5FREA
QmpFOJGUu5fbc+qGhhIY3g1OFRWyBxZuIlafi4ITxRR5OzUfr2g/craCvul+s/xnvVPIEzxSPHWN
nzONd71TmMOxUec/meVwB/SU8dPX9XFdsL2zb4zqmpTqDaiTqYuU9U/i9t3doEoA/diQWx6LRJdd
0HXtewq7ErnnMht09NQ8iKzkSFb07fR2ou9oD3Q/9BfklT335osjb3A4aMin1bkD7glmgAT6nYGH
sEN//YlcoBeQDo1E5sejtFsCcBk8p9u4iLQXn3ZpsANRA1nxkyYwYjGM+gdYBJz+fLMcU+qkDWzX
BJPQYypPeDQAV6uviHPzdMYs0lGjNbUnuXn47II7/2YPqksedTBK6fl6f4NrHIbsbNjIErnm09Pb
MS8k+58poXM+GZrov1FSKpyCaym9w/Ez8wOQG/fGMAjCiFZxrvKOjyf6M6P/CMlp+a9mKsVGDUud
a2vsh9kyrXhEe8PCoYgHCHC1Czpv7RKNbwXlLiL9CmXvCuyQd9Q77QWdC52DA561ZgGmHOF2E2RL
9ACIvF/9NrB6ehDMpwMprDRiuGJ9yMy2Zcwu+tP7qwdUGcoGCAoJOtE9aS6dVlxc+n4vP8NWIE5r
Cf/xw8py0ygevopPIpPjXZOHKdsmVAujuhY/TlYDWvdUfAuggKGY8/jeAJjEUvYOgFqFcvADzdd+
Uee2uR61epZFYNq/vIjSKzRFlDG8VfXYDhQB/sq0HcXu0aPhLatbWrkFTdztjfTQ6JugjPF2B8vM
J+2lEHsGJ7kfVrWgZNjhR2LIUMSf4L4kZSOtkdXph1LvxK2Z0VaO82unFaSjOWK73VGPzYeAwc1m
ed/vVh7aBGveYcNq420DBjWEPqyRl8OK6kmI43TVmzyt4Z21JvmNneQevqEVyKCYYagZieMRJ5jT
9ta+QHAO5Db7E2CjfW8+pwc6cFruAMKeyj4n351E90BUVrVqPB/eVud99LkLHjVRLWbN2L5Eg75O
YB8P7C7NswiD0CkLa0LXhIgEFHDMaoNs6z2j4S6WOdMM2q5TCeNSh29UWFp/hEv2DtYOF8743LK1
YzWjaAo558+XGZPNIyOwwFSjuocJrPDax7DulaNLcXwC/tO3DPDUPuxuIu1Vh/2ty3GPgcLVxDLT
Ek4s1+Rt1lsvjDJQOiOFZXCE2KjrG3+M/ZwHeibLtdHhznQHhK/vixwJtAtLhWvGiPTschqtu7TV
s6A/pPGnNY9froYc4ZGnFVZf7+kpFmczP9mS5PMqzpRXkelfZOVGatlaYik6Vs7orlsy912v5bhv
YfhvCA+OpTloL9b3QnXcxszdxHCoWiz9/5OnhkVqNEpqp2aV62bywNMW7F7n4On9hid5AeeBG6xx
HzMH5EDtMYYBgY/IiCNsB/ng8xuIHzVBjaScVs1sOqimj5vchXze6gth3DUxUo6lhq3QPd4aZi7X
fxZJSWBq+YYgDzLh0X+8+XSEjZcST7gZ8BkXlnutwT6aiVDqw0LoeUiw3YnykshWu9nt1MhEA6Hg
NmAY+q2/HgMTc30OyAKE3h5VN5NRs9z7EMEvdPViUnptU1z/j1b/nmb6y+jh1ZuoxZZCOQZuk5Cs
T+uJa1CSn5yfMDexd5KCIJUePGlWmcTR+JiVPw+wM/08L6vr8mEDuuTG3AZDoGmDpOYzJ9Z1xdnm
PMsQXt9B1RHPYVdWTnK62f6h/zwmzAQpZG1Z0f9eJ7jINuuAX23tyg/mFyLmCgqXqEvwYPmNiqdm
3x8ZXWoUjbdFdoogRUFgYSp4QhWpOTP+Gn5ztjCE338I8YutcyghBumLmrCEov3AeJccwJv6LlfY
b5spSBqbPMPsnn7OTdP2dTyRdB1bufrZN0Mj47lnd+4VVOQ4CzaUdMGGDMYLEml23GhrwM62h2uT
4C2De9xvfTtPm5StkPYTP/doR6WwSAkvLpnW6cKrJghg+6r2/qxVWix7+DcOE/uw/j9O0AFp3olh
TuPTwIPb9iLGwCH/U9rW9rlG8ohFSchmuScJvwzFBVZL37+9sHN+cVeq1qlKdjp48Nbb5dlje/yi
4Y70mx9cq1bmz67EtpJxj40NAlAW4c2NnvuJmOPQPmN6uxXIRE+X/9OC3dXxJXYfEMAJnKQvilr8
tbEBcrdFdsX7McMSVHkPEG9yNQH0liV9C8zdFGfFkxHqYyPbBc6MpLyq53QXUwFVQrx8F8CcDjIB
VagYQjtR1oLX23cDakT/pxbNLrS/pXAT08Zrg63ZzPxcmOPHYg5oonP+7UTzxYMktw6otCuNgWT2
M3zDpuNzOZ/vWoMis7t9/FKNjB8nxuCFrNV/yiO07p8ezrXteVeOcCzlG8xlOhFy+GY9AA68Esha
CFw12tAk7oUb5KAsJFPfr1vo1Y8mUFyr5l7cC98IUitZgFSXVwC+CG/0EFZMlI/D9EEfwGCoY1UW
nrxE4bpAYhG7DR7dSgAIGQxCJag6OlMqQpAFuHFqUDs0so0euGvo2UN8XFXLyt4QUMAFfrinjltX
CGfemfX9VjdzuDfBM6uSamhUgYcd9OyNprUdISZxBR16lAFIJ2M0xYLOTbWH1j00I6C526augYrz
6X3mVcgIvGSb7rEXficPp/IXicloBddalLrr9O9N0XYnfx56vH3x3GP2+DkaUskO6KSm793F+0F4
b2Tq1YbVv1vp5SJzWaFMq+A2mLqO6Sq5cbCpPFMgNb8gAasw7n8iZT9ybBF/MmKf0OUcayhMF16j
P12bJfIMgkzVYW/9iJ/hsWXUVT/qA0n2B8MAAKCeaHvpc0EFx49Y5AhNwupNUro1suOdEtsBEmnI
uhCbihDJGk5gjlMeeN7d4nP4wmxkZfovyzaMK2E7HvGFl3OuX5PV1hpxUk+VWJ+UQUNlsTdvANiy
L4eujYAKyjT9X+tipOKf5if/GWwqMZp+zJefGXDG2WiBTzhF2OaPLXhtQ3VSS2/8QW2AIi3yQg//
Mo8DR5Dr27AfmTqkxtXZvw1/0qLi7yT39/HQKWI9eQGg2q+lSZXbVqGFpwS++zWOIWnASo2J56mB
PRK62GPp5tzIs8vbaAZxjjh17170HiaOVra2Ubuu2+EoIGMd1IpdTJt2cgmLrKSr+97+ctpl+vGe
+fo2sa+/pO9BFCJ8a7gV8UjbCxDYv7wlbUOL/BUXJTd6sHZq+oK18GruYhOglgwQfzxAHcEN5NzV
3G0U43xoYlHk25b9TRRZBCE//LOS080kUNGefmrFdzzHXq20bWnaFHHXvUWGq59sdG8hlqFNbDyt
Ct6OFET0a2uU5ONjSWEk9yplBng6wNsSs66fFM5PFxgQNJ6cc0w9efYxaEchGBYlzE5+0OklYuoH
3+kgJ7LYfuYAL3TGSV5O9ctOzYKxCQ3tnCRJIDasL5u+W+3gj3WHVIx2J+0uOTecUnCMPVLnfAeV
wku3KFalg92cpQn0y9zUav1TGaNS79CtaldCNHNdwStq5usboPqnJ6qp5agvfUjXE6I8SkDOSeL6
wdkY8ynRh2F2vohC25fgtSzTUYkNaI/iER3t2VjkZcwlKbNakD4VQBFrkBzdI3F7fgkKsAtlI20J
nPo6yvoF6TIesABPL25l6gxq0CkYSjeiYvVOw7MND8OvNz7PPgWwVaywf08NAoeihMy1+XEJR61k
k5QW7NFYqV+iEf9rMiVTnVr+3seSOksRpD3axDwCHLgYx4DmaXvFflD8/UOJZiahGl5SVt/CbcHF
yEQ3fFWExslS+wxuOCriBCjuvd7buBxjJNEMaeJnWb5ZV+F+EKt8+bxFrRsGE+CG3d0LkdsilZnB
EkvMTQ3ONJMlwYfnI4WA8cyHcxubQAQyFgO5+FvHpLECjds+kcbdyPeYKr5pAuOMHZJ3J5mBgQyH
UOiR2KKi6tHw0wFTpr1L3AQLFL+cATNtJdwND5/JduXWP9+IyWy3Q/W5h0XvuvhzVzIxWcdl0zG/
PRbrH3xR0larN396FaDauVUGOj6eOtJ4s7E9mdH+/I4hqZ8UlvgxNAP8hC99BjhCB1d2M3nR3rtj
wFnonrv1nXBn2gJke+D42CXZktMnEahW0888HGOmfKTnCDRKXdBR37DQCyW/gjppT/Ha1+US8MdA
ZL8Q5t+7DOx2uVmscWbBSHwHfgEj6/4H4yzyz1lGHZ6cgiJHCDaUTIOFXs3YrLcX6z6HQAwJP25i
jzG2K/MhEvgCPFxPx/XAwau+h9Qz2IskHb4aA0vnwn3dqEzohT3TcHf7GHL0mWpUuoYpKpwCT/Rn
nmwtr5qtRIkLMcq3lfUvnmRYoXViqmeR/GyVayPxZxouA2lVo/AnoUP63CaiVdJj8Kt0WByyjMcg
kst09EVIy419gMOG6hJRyoyTFAwCHRS/JVuakx+T4vQtabXOjy9vcQ+B+j8fBdnpXVjZT0NFCMLU
dG8QWni/I/PulI1KHZ+VFw6mLSgIERy4tRVIMkSZ4wNim2AjGGGzMwDLRStpto0BvZQ2PKId2e9W
8xZgth2KP5zcMuPTLrpd74FvGRln2TCfokpCjobLmoRExTpJ32yUr4DGVeIWcMZjdMAEDUGgoi4e
UrEXNJqhmTknHCBWd5c26nUdVnJIC3ufGsQphsNcnVrTuWI5g15sLTrsVak9LDdmbnu9XLnm/P/P
h3LvmZ3BUwrYWLtbdF2VF2wvhCWXEVMIJLFVjb1Z4prZuNm/OjmXHYjRThTmOKTWRyhBLwwlXRa+
93Psi+p3yBGote+WMb0cj+jPYMm9pSrOQc+xYUmAhfj8OSn2nHRJ/lh8+BrLC9UQ/GxuM576EXZS
dv9ne3fmdUtGyqwlas9vMr1jkoQa6cOw/gMxxkOx5Di8Fsrpvv0iq2QyOpxcD5AQS283gDB90938
uevlLGx39iIa70PHdWp/S99XEg/uYYZvfw2+bLNFdrVdk+5k31vccaSF/F7rrWAU6AW820mCz/kA
tA9rOSroyGKhm93wiUMxw3E7bfYwQgwR8Q9vArE8383aAYsfclmF8bF9iPke2KXwFEkGNXHyUwEN
5yfyTgyG2fL0+i5YrfmjNnyFFBDdrhZMn16QGQIloN8MYOSr9haufE4F2ACDsXF385bwl9bLwcXL
SHl7FweXijwWIHOkGA0ck2+wu8LwrTNEXr26p+imPXUagXMBrKNERRb7/NaR8gZGr4QPFgMuEnMJ
/rK701s37QhUjfJUj5wSyt/eTKMbieFqRnG7TdZ2RoI2lUxKZJEgCO9r1bnGWtxaya2/p0nOeA3k
j4woo7sHmKskmj2Hy7XQPMnCYj0u/snNE+0dzb7tOSBhHmA+4DSJbV1qJNrCbCrY28V6qiMStE03
5hIenLlf8UDKsPS/DdlotMjL6x5zY+azGwgr1Ym1j1MdM3TNtneH145dpdrK5frfzMb/+Sbhf5v9
8tTZ/TckUw29OEHUFiPeud+FTBaYH9BM2vluwhlNKH4B6Le1Podv44axiLvcerdr+magr2w5NKd6
zvbhTRTgDigATI13aayrr/iQE6eJXJcTxPUH7ZpjOlwLQXr5y7/esotY4cd09qPsYpjY3XY1FneH
vabVCsjtWRqWsmbN36YulDE73X1mBFD8xVgiehptFzCO5ghQohYxnieHPo4NtB9xayP94EgTL79+
5vUzLD1l1cDrjQHp9ysd42FkgRoHBCGy0xh3avj6NmOgTJHRqxueVQIkeBb9qLRYISt/PvFHsVtD
QXXCfeWXJ2ZTT3joj1MIKeHhOl/qpSzOhDKnieZtTSYBdFXEKmFbhQnk9er3WVvx+tBDYXJDjlph
bBBXiT2BTiTwaoIWClqoZtagDZEqCwRR3yjk/hEcRO8cxicG9UjoQB7xMocLORA7K0LO2uC8xReS
P+qXWzMxFrleQ8fEoXX01yux6RrfvIzUaBHcCcyBnJpOaTzYVtrFu4Cuq0rzIZhKnTeOCnzi/1we
AEeXI0bDBN17E3x2bK9wIWkgzddG+l7sY8a739UmfHbnPl+96tzSujIeAXHGSathczoPCBaW6f0t
HsEgfewsQqr/GDGv/VMh+1SKJmsj9t1CgkvmjsVQFoT2ap6iaAg/AdYx0iS9jmcAchNzgZx7ixPy
eGE7TNFAhF3G0KBT1kOvPT4b1hp8WwCBBvemC7Wr4/WoscYsuJIb1J3CXdfJa1iG4RV0Kk3ZnV25
frEPctwDpbUpa1lPAXn/3Zn4V2s9iuWKYO2tkkAWbXLUlTQ0GMO5vNwZi0WCgX9nxOzuSXIbA/ap
rjjJ9wmqVNMhwPNpHzBTUoD/GDSQRN99t2ZXk/M1skaX4TVnmyRM1xwJu6gyFsY248wS8nyu2dvi
CuLxvBBCNUcqRFKi8d1qINVyxqVyj9qzlY3dpv5mVU14c/YhFPmZC/INsPhyNVRvMzoQPdfxhh35
zPwHw7xFsG6lONDoaOy7fiwMhkNnK6d1ZFemwjiYsqrMhd0/zwlYYUftDHIldlJhoNehSe7b2VKj
heYpwutrXOM6xIW5Ypj8F+Mz+hSnJdw+uPkPoy8B1ap8BcM7eBy0kfdn3ktjkWeIyhweLvKTpRWn
gouJ5VydrDiYQQNG4loVD/U/9fpey5rSJy7fFOxLsfbXNisUAfGCHLr6ieYhy8qcdemblSH3tGhv
Arlfub9juZm1UzvtU8MzU7rWJPKq8/CzbACSrnzaJkUf2/WUctzeunUCRv7RM0zoU/nYu2AiNyvO
yU3jQi8hqyC9R59HnaFB7V/vIhsGNSFIyaSxAEngy8AcIkKq9QR6eyrapAVZ06QJBrsbQ457jhH9
GkTg3um1HwUHOmFcGDnxK5uXgLLwozw6bzGA7gVl/J2g0CogItJbm9fVdQwVSk1+J7vwLqa28f7s
YFA8ftegM4MxIXJf4RhHbLuBP4QXYlnzrHgsN8DRR+uN2p7rogZR/F0INr/i3PgMjsG4Bof4NjJV
W/l6GZw6nJ2uko+Zh4D2xYYbu2oqbLPcbFXj00BPttC13DlR5jpvvasr5gsV7QKnyfdWwFkoC47w
6rJQfl8q6tjYLn0Z+f/8pLxE3nf7u6Br6oeXbxRM5JeRJrTQz0QuDzwbHoVT+zHvhK/a2/ncg8x+
iLHtIAnUEHkrMXX0meJzhTsfGkxtVMSGjHsnT2pa+8TiExRKE8N3qMWXUYHRBCFt82Fkq19TvhGl
tgfJc/Hsl5LTbrq+K9GiTc/MlgU+n7tvuZu1iAxh7y6tJfGx91C+KCrUFgpjY2C5SEn7HKM0lPyx
tUgJr9tet0vaXxvfIW23paEOWzoS3OrhAHzbDzHHCEqTN4p+9MPnLzD+tORY60F9L2XfPAXhIFTH
Q9z99bcmYWbOhKauasfMEF6nhfhH0yjgqPVuulhxOujGj6H2d0UQV+tgl9HT+Tg9dSYJQ9h++d0P
/vROsudJTi98vJVF+x4thI8kFpPuvkgaG26D+6ZAiFkHjTMryVigWCp0SYWDrSxTRvgc1gBUYVQF
QoC41wFh+niXdogkSFqKp9phw2mj8XQT7C8eQTH5BUniRsIHxjOJgd4onpOpmPPp4QBGs9XWnPJV
D0dPMH+km80+xN3Q51dTjihQpDIVbxp3U2FvnBeaJq4cvNVei0TqCgTHah2V77k75sDFuiM6Tjwa
qxXBcS6DvhUJaIUEEparXdqNr6AfPhE4q3nqr5Yikk9VWPMhvGiVqr7r9sHlBf0NFa+yo5+U57GS
ohX7KGWo4rCi0NXOPNaCvVu+lbasV4wKnWyirVwkIyuXQqKOO7NNKVC3nhcq6/3Zt1sMJbKmZ2R9
1GXmANrE+dQmJgXZme1jvGqVZqxUiRtkBX6R1xb3AMxc0Uc+K7o+A8rw/uLX+wice0USqD2EYNZ2
ONboBBPxRhzm8efOj9ZrBeYiJJU3KmKhi5OPRATavqipOO4HttuwOk76FtKBwNEo/crMCZwgDV0L
Txtn7ik+LJnEPFfH4soexTf1VYwZHLb/psClzz47an/643TeTpIuhHTii9sF56XFUoVkBnRw9+Ff
cyEUCTqLDypGT9cDysCMGt9At39Nh53DYfchdFMQ9QMW57iXmp038SIj+adXM7sfvDp5LQP2/Y+G
gompKk6qvyMiCZ13Fj75uBPFgBOdPyQxUmqkzZbTu5zffYLaPoPrJiMn2kyCYmpDFJtvbCsAxhCz
mccn3YotSs2tXeCog0f7UvQd94eyyEbzw+AbNMg9M6u5niXUT+2i1A5zmLdnjjqWxJkQtElNq5gv
mnFxo/pRRtzSpPsfOzmR+3FVb4GvlvVYPutidzaOSQlQS9MO4vyKt9tLmnr1JMg4gCSz7oVa1gUb
hl1QMd57N6rksKI4fRj10Ir6LHZ93IdR26F9xFSRVmut9/qp+xyTSh7t2N2PxrJRBiJ/seF06saN
Te52MF2M7nsb6giL4M0LlVMOjJBwhS5m9sDmb3PSV3ZThlhyZhP0KM10uyygPm1LKZNgq2/3yIFe
fLRrdgn/wZMy/bluK6D738reaIX1UGhduA24sjIDaB4/ylzQcdHZ1N/31GOO4b8KnQchMAkcxmAO
IiC1mjhGbF4dux5oVg3CRRjfOjHUKjLVCbVgjzPKFLXIH/WWjnCVD+9PXpb22lenL1atKjBBi7jn
L37FuXQTt/dZJkwgBK4w+8Xba4opZyUrAO7dPu8YFCI4SW4aJbmsBmqGWEt+HXbYXFqyqR9ucwsd
oa8HVDKV9xOHBSoIlfVJejKUs1+NtzpC+IUgeg4w+y2SkbyyD+aPKvJ/hBbxVby5K3u3Pwz4v+ck
UwamzGl7xquMm10MR9MSBsY7MQLoY13xniJ3ktAY66D/ecT8IL3AZz70kYzst51ltfz51tHMKRZn
xgUEgj4x+wHW0ktLkm8RUOkbPppJBWANX9sohczyOUgbX52w3xqk7WGymk6nQZefXZHT33ydSS8E
geCL2M2fMMDQTc/6P8zVhm73xJ3m4QUqjVO9sTXxbQhGcQxeCHcWqh26ukNVbJOHYglsBF4P7YQe
lXbYHRp90X4Ba5f2Epyk8m1Jq/qAdqWmpT1F+5J4MvokzjX55pwICnYrDs1dOkOPp8YB2bVmt6Xi
GHzDHoFyzobvZc6YSnQAx7d+RKyjPbSfypnVWYNuTeU+S6YamvFrb6OIvLmWvHnHxYUMpadXNgl/
mPcmAj26upzii0GJ0tEkSLwQ7AXJHzKbUiFAuKokXzggVMHVAOUbh+JvWJS2O7aX1DOne/60NhTM
b/eZG1ZQSkfcFch+4UOIfsb3+60JLagGJ+jwPQOiPoMWrS4jD005JYl19MSLuFSgjjsmfVAKFsO7
SB0sfE+tsJ6JjsKjH/WfN02JC5k7jwmAbfSzRGbu1EBa9wCuk5UjwyV96ardD7cSpiNkeCcMtb1w
uWF1h2UoHlmHCSEnTRBAI0e5VuWUCZobUGMA8FqnPESpOtFSAbYUJmGAXeoWC+sUWYJHBN3OSwuH
//1ersz2R2XkAhxWiAYTm5lJbyHb6DFwcqcZ5FJarIGclCG2eMckkmlxrEcH8hx6A9QueHeW2Oye
xSoxasnFouqwy3HFq14AbdB9YrDvo1Ir5eltNI17UgT0PYX6NCPbgy/L4LGI9N7wNmP2N93SCOF0
99+oKZdfilhCkg25qDH83n4faI/rubu1rC95v74l2cRMKPO9eBkjk37H8MxPrn8Yep29cI2Mc9ec
PFZI5C9aBkCqG5gUlSijT09Iw5QyI/afblGeIpcIrPJrJs9sCPItox0T7kKvvq0vr2a3NknQA1Ze
l3DrZZugGVowqg/TG4sjaxDY12H4SdCnEhJBEyXfhgOPWozu9uNy4BjOqy3P85xM2omqVb+oQbdw
HLqjnqRBjLiss3mH65NbEeQvyU0RxAHUlE41FZFDc7un8wRF/RahKTDdCWCWBl96YaY6kYovHNXh
pJ51ACM7pQZBxGpysUAtyWg0ZYgYz9u2z6WxAyYZnlAyzNu6Vt+03fmLYOMsINXeW6XByY/ciIxg
j2eGx4oDBmL0vYJ0+espUM4XgOmA32jiEZsgfjjq1AztJuEupKhzBbjPpmD91U+c/B7eQgGIpofQ
PsbF43gW480tCvq7C6yAR1EJFzsFnAj+pCkiyTSm26rKMoJOjXDQVhUhSxG1G3HZSKNbVwDGJdcM
YO700VknT9js7j4/gakacaqp6aP1Qh+0LKD6l8uXtyyhtIHUXB+wigOoow6EPm8eVslwjXW0dYE9
3NRCnnav/SKQWLcSzmauhOkzUSF4hIw4z+WYBl/b05QnTPq3lYmb+tE5EmKxp0cnqjDlSGllPYzv
x/73vhgESJt5LycP1dXx4dWVGAUhG8XmQ37QF8bzCfFTQK1chuZUyE48hdDKR6MPxDBeESvJIH9t
3D1IELVzD3Poq7zUE/HZDJDo31TvNV2WSzosdsGj1IKC7Rc2Ry9ATxd31XAy536J1qmjPu21KZd9
V6g6cqCG10N4XC8leTaiRJHfA27M/K+pEtZj2qiZaZDs7XDIEAY4lK+02oJs6MKeLGV827/ub/VT
/CTagaGUuJKUydX8JqEPIgF2/ShinfMLBJ2i3RsWELVxNyaB6Qu6CT6K2sNwdQIm93dYwTXrjQUm
HU/MKH7JJUgvQKLltasFe07/8jmrvRQ9SCNHB/vPZIEKWoz/Zbzfw3zinAR9uAQpBWn89IUw8LlC
ViyQj/5wmQ9qZCw8gXYFBcasKLpbon/S86rZlmiTCiwh8re+yoypVhKs3qsNhU5XQJZ65iALSJhU
Wkr+j4HG6avDRl6fcMVkbqDlhDZHql2PfiGu+PY6aOTso1hj9tZNlUliZn+V9FN3Y2HtybJhy/5a
+6jRXZ976BHj5jaDAAe96msr3dIMBfJbzWUHfbHOUip0x2/EjssAWAAwSwQW4oG6+eRm9c2Ki0Rv
qmKqBcYlRgBVX0s8hT79mh6i2WMlbCZg93u4iDbgNJjQKgEnjxvTXXCO/QJloAyXi/fpW8xuA06X
lHaug5ox1m0ngY+TZniYI5u9mwtszbKuqg6rqt1xK/ADxyYuiJ3MJHsQtF8kWnq/xE32Jcf1raPB
4gBsWKyAQveJk2ywU/bIMKuEMMhXhDu+Mw/QzRNV1hEj5PskJZqKyb0amRs78PNrvjeZmypD/uUK
jNPJLRAuks/RYndi1PQEl/atEENZCgf/VadSOTklPycyniAqhqB6pymwx2c8qOfR+TokxQuPdJ/X
tEfpbFoO0B2YL3INv27p451wc1rArIxlaLuXoXipolk5ng9XeyMTPHZDHBQsOOlweqeZtmOpA/SU
Wdm/+oTrY4Qn56+CW6E5mMhIPhWxDEnW0kD0lL7eiup88qUpQosSgBMyuE4G8KbjTBptHyg/e75g
8cYUFIcBEVbbcTtgxdy/Q1Bg9crsjg/9uWiqqmcZ5H5ycuxWxU5LUaYkFg1KcNHaySJtkht0qXbe
x1Bh1b90/SBELb/leVZFNdjkytndxh4538wSvEWwhFO6ZGzMqk4eJbJW7BUonEITYHb3Fl0senIR
JjRG+vEQar1FOpPt7XCndH9j+4dD6hVotlCOMbznr0SmZB9WMLmgn4t69soIcfSzs50vKHVV6+Bd
AE3Sjzhsg9zBXrWymnPT8wijrOkFZelsLe8uVk+sSvJFQg1vTctVRBHQEuiP9FbiBuXNaZi1dWG+
YVjwnV89jbk8/0hYnhTR88U4rezNMbecR5QQv0hYB2cKtdnZMvLeo+h8xEuoK6j7XpS3zqSCCqfl
p+7WG9MyyqtNEo+FUKok9qFfHNILgYnfjs5qrcle7xHyazEFqLmkOIYOFAq+XgRFKOHS6eVODTPT
CARJp5MRbordGIHlsO3MDfG1Tz3RDcZL732KKS+Dc6y76U4WTDbbu9IzyAtvg+xd3ISrvF00LNXx
SkiJdbsw3l/x7kP+dL1ylt/rHWoxM9r3unYH2GPKl21PYvusX/ZDAj7lJ8YtEF5N16Bj101vWPda
6vYinv/aISPHYhyhv5UPXy3JN8fTeSy6G4rpnD4JFxBc2XmmpPRI7erGwzHjhsZ76Flq9nK5DPXm
O0j66v5Zbz2jQmhbHnLbgoHlzAC2JePy1+P73u7ielp/QyUbnRu8U3bYCxI7d4JDYv7vtQsjti5m
e7D3GCunJPcsFeud14EZ2fUVkZiTPja7h8iYVRfWZSwNWwVNbUkqkaDlFHUGsljBhX5mCHOAJFUU
aGpblmq7nvoM4oARgKswLaZSYKSGa2JTnsoOhOAIzMZCuhYwZSkgmb3kZCqaTa4zZquMMiglw5sT
5CCCXWfxzj6oRIYl87N4jEQ6DpYZUeC23rYtCbJBHxE+kfZvle9dqSewaz5GWVldrlufat9rHpTg
FWBf1hADl1VPr5nKnYBYT0l1naTJyIEpaoGboYEWhRZwkjpGib3GJJH1qH9AifWwTXGkoB0wmsvL
fL8ZgEoQDyLQnbdFM+KsgAt60k0wHYuoU4ql4MNTqjY5G1xTLJEf+14mQWRDzPcPh7hPS+4WsZb+
jbL3golXj2Orw6ppzrL/8LfHAonZJ8lEygRzeqRufIAaRWdfjny7rSMo8jRPatw7sYOMnnJysLYu
5zXX0vB9lpfZZT0tb+hOI88Qiy+ZxQZ55TROMIUoGK6x+jauhsE4CYBK+wImwXSVjVZK05THqB+L
mLAeeyD7l0CYAr99A89MeuiZmaUl2QPud1vrQJ+ZvPcX86qtXhijAwhIxzCFJBzbzIDYeDIYvokS
4az1Ks/9ZzVkmsBNsOM4rlflAoKBs73pQkVHkMJKBTulZ/X1u5eY2q1esCQfur/k6XAJfTi2z3Q+
tTNpah9eQ7f9wDZKPhJgTC2ET1AiiS9qCsnf2EB+UASYPnIxJVP0apYtQ5Ecm+YZPNe40LeyTHpV
4fJE67vwXESH9VVdCssdqaDkiJnA035q1Hf5eBblfRtj6m9to9pw4JneYsblAa9XlcTv7yj/4yaN
XROfX9lxR2DcACW9+3ZFxXOHq/gnOuG6jyHIuIgRS3O0Pp7LCOpDg+jd7y4mqnchiH4Eg/626qm+
+W2NFAnpeTPawPCoE3yWWk5QUk5PAUU6EjfowhJlqpzWm6hzjjkklS9z43/32/ldLSvoLFx86jha
TURtq3Y0WaqwaZAj0ygxkctQgfCaV9RaNDeN32ZCNA1dP3LgnXBQ5T6ISqdoGvPk+TRusOj0+dwy
18JNDNa5FaIwkUJAkWZ4lCgqJEx9ExXWso4PV6mSYE7HWRlFvy0Kti7TMWwEccWXksLpjAmYa1LT
REhqVbnOSVxURvBYVOvltBuS5wzrQUko3b5sovE4j9hP3/bbwF/Ge4EDKG/o2UoOURQPG3k3WYcI
XYUNnqSwnH7pwQFCE/wHh79MvMci4n4jo8FtBUZFJHEA1ArKEi4Dvh3nLbU5Z0ALq7+Qk+NT6xbc
IKvEoyGNu9gyV396soxiPvtygB8p3kR4VAuy+/Gj1JKXQtgXvIa99KAl4DgfN6OPCPCHKLU6jvHn
9yG+2MlfMABKZOnAw87Z6cenO2ydHzmHmFQgKFX1iIZrF//lOSqtuQdmKjCE4HazpRxNzE4dJRM/
APzRvf3z98aJJod6XusgPYvMqjtmfOBQWI9T8mVa4bOMU50TfZduDW/DjlizvhHmer/TCtZMyih8
dRvcLOVasrEx6zUbPaQSplhjsPNE2vmgJrG5dxqGl5fQD/SkT0l7LrUw+bzuhkZNYMw1MwNq6Xx/
17phcpKpt3cYorWF4S+7RMJaXeTR54fUUgmcn69pShBVQsm7n/oMIFt6//9psftQTJJB+hDcbUda
dF8Vgmrroi3UAUTMDIAtkYwighHgKMT+/jBVFYtNHeFSEUxd0qjsDul2WdhhqERoPGCNCjbWWU41
3aHGBkH0WFRow1Vy6CXg+hyJJIy5G+I4FaMiQNrbfENHk6yNWXF3lroBjvuUo7HYJfU4MGJ/c0II
aQGml5e1mzIiKRk1TaL5NqKt0icKRsIJQIeMMu7cG8fl3Nj0CmHOAiNv5C55czGFv53TBJD94As7
qX/LaHInkKqYBJ9tZxRYApSo+aEoGE/BW4YS+TRmAYYr629dcEOqCBGBmgrGSNx59788ypoKJptD
4d56UuVbRZ4zaZH3L5eSlUQLs2Zo4Mt4KoXVktz/LmjB4skL0k8z+MZ0wKFQmeUlKNsZPbf5S2kF
tJp+OslfyKDeURZwuWCxQ2DWeXsbr7X5UcxtOE/GH/CtGeUw0Ar053lyzS8SCTx0DNtEN1ojvsE6
ywsK+6UCSSRfQolCaeVoztW5vpTBGcm9pGysp+XM5T6/brU2ygyeYObFBsO6qP76s4OcqchxOk9F
zv1g5/43H0tZIFTn2Oo8Vhj2j1EbTZO7lFtAeWluyxjV7XVEqCWagMVLvNHvQi8RWbS5ATDJDyVu
hafDrvaXKUlxHr0jrjRvVd5TAEgWhI91hWyfb4DaLdjbO34sLyRJvK0v+4IRalGmRdhTM8y6AuaL
01s5W85XTz56Q6ij0L0WcsKmvyckybRvmr9nBpoe3FZA7n8wB+ECAH26R6KkYhyaIRiH1kAqr9/V
Om6Jed0pyWtg2E/rm0uLiD2gMqjPu98A6jvEAZuBVillwOEt4q9OSmjznG9tEoyaIYgtXmU+HDG/
cf5cDHWpR6qI2DNczf2MF++2/kuznbNnTTIrKvz7FAIcS9gvNRJKjT3CnnX440uKqBsAeXJipAED
M61UZEpjWC1+c6+293R4z54Ok1noniJDk5NueVMygbUMEvM9sYTZNjc/nXAIO/0sBq14LLmzlHWC
vsgH5ddwYi/Sp3gwGeyV/M5H8OwJP1CDsllWR48WNA8cG5GnNZZEQ3AnHNmwODmCdD51ZmDsu0Oc
6DREX/tTKdKtn6bOmRDUz/WbSG0ut3bmwucVdzIR6gX+ARvfolzb6lkSuAC7YTX8GdbFXBJX9diQ
1zXu5pNjgTzjuvtu+la+86lpmGaa9Vd5OB5enyFlnupHubMB6gDKcrs5TGN7LEBLCIgjNb0lHYMk
LacU207D8jnRnXhamMEyN8RqEqlSBrpgu17cOF0e1IggQP7LUeacJTpVak/y9PYqxWsJohpv0/m2
pU7LCo37WeAhGgkkN71GgfDIdCi8MvJuXK6Pv2nvGbL/P1khTCCKrBRviSEMfxK8LP0Ubpwnj1ql
sBs1zv82KpGvJl6vMf76tOLV+HgbIvS4IvlJMrrO8DiihYMZGccZkd5xgm8yLbJEPLRR8OurPlOR
g/9tIuZ7+Kg2QpPR/3uRU6A6g6psYOdo75HurEDeRWzsmXPd2JpilcYZa/OC6IeJcp1AnvIFmjeX
8AZla4NV91oUcQJsZ/duYitMtK8X1h+kKC8D9sj9iYv15BdEHdNzTu8Gq8EG+/XMR4Ql5jx1UEFm
KVnNPsL235UtjfV0ljtDPvJPg0R6lF2ap7scvEl+OwwXLH6JDcSW2vwSSnA29GGMEH8sadeCpQyB
jnmPAM2P/kdsVd/aRMH2gbDzXMkicbb1+b4vDCcHguAF+XWUNJGP7WPQD6X6dZ8pVnT6hxle1xLH
P7bDwiJt0B4J5XYPej1Qhc8MVI0BseCTHlHi/1V5Et+mIvQUWf79LeRMUvhwTT1HeOvHD9niZ97u
E3SwTleF9RrsrGP0G5f/oN8u1fReD6SmjpL2bL1cUFOCESSDXUCwmDRndbS4BX8teCTZja2rWIat
NYmui8yS6R2GtMH6R/PohLVfvzOovW9gvqsRuXk32/7S4/hlhAe73JUZMwQ7zN7gdwvu6cf5u+Vz
r8nWmTBOXFNuk7meqmbh8mTkaJN4AHMR7j8vyulFeIME/luqi8hcE0UKzhKaXwruJXLvxBIoCL2j
l+JqZBlDaCgl/qr9P2mnzejIx+UiI6kdYJf9SVdOx2vIYC3rWzQ6Z3xoMbIt28QQIhwg5hMZ+QAj
5Jf+9BruO3eVN/FUSwdnBHHHPL6W2zFly3MXQGqJHcIoty+KWj7o/b4k6utY1hIa4tkSsMHk+Wvl
31wElFhY/V0oLZfO5JEohXnQtfubOn7kRkRH4YaFIduYG1AoHwQrJu9OkXNnY/gapSibmzJtrpv4
vxzdN+0lFilqxwfD5IFNfYbFdpX5fiz9jVoqljc95BWUR3Ywe6oL7l2HYnbYxkeSvc8n6VNiC8Uu
BeYO2PHgIUwyNEJfZHZ5SHkdmq+e8Z5uRN0Mn/fOnhkGzetUaIobaHfx3zW/UsU+Fza11fGz93Je
dVB02xtjFo5sh6e2aL07qRmtFdQQfJtLncNoumYfjl9xtu3eW0BKmCXMqvLb+KGJx2DnnIcxrAxd
df3zPUXUiplUrp3HTx2GHh9fjj8tARDf3mNX7lmFlkus2UnbrHYktegshVctwAexXasx1NgDuqWf
pzQwZRYSk78LA/oqaO376KK4WZWni/KX2SJEMGPuEuAK0UC82p6Qn8BxoTfxBMDfiUQ4bE0L3Bf0
4yF5lHKT8sdU40Af9kMmYqVCbpSa/isk0vNtVb31I+cTJe8DpDiI6HBrjoHmS1cbPKGPPt6lhrgx
fWSsfYC6Bnxw1kt+6MTGiMlQxV86b5H13FGh8FqZV1/5jstpJuYO2RrBkqYp6VeZmOF2DoLdT0p+
A2pp2ULbEsUxgumKW0olUqDE/t3+hUOMaoEQZba6gxu9Y9YEiIIhOMVnpPMCRpk3thtOgLYxKQ9d
xAaJ9MvUIeP/4VgFv74W0f+ZE6b8L+QGnJ6QUIzQjXcSzOmAi75XdqTBXvEAQl+q8KFJwqg7pds8
jYEgdSw9yXe5Swd8OsirZDGfxAn1ZSdDyaKOK3yIPNXeejv/7QKto+enltpvk0yciE4SE2JkLtnL
uUDJnAs5EPze1aa/l5TdG7cJudSNwwVrDdzBG5oV/qaJGsvpCI5nyRu2kX43XD1dJLbL2EO9eKoA
UojNEC5ETNdkyuVnU5/Edk6+4wyyORX11hNfd/0NAl3AAgp1rKGV4VqF/u/Dlzd6h57wkHfwDXJo
y3FqivT/X2LtyNUrbF3dRC/1yEIH1AtDbNBpNP+XcBbzBZk50Z4Uai93PZ/yJJVbwEK7JvnxzkPq
x9dmuOSfXaaBwPH5fnYwJ4+48jygGMNv6UIBWTTRQ/NR3otBYk+zVUSm4iF/9TsbbS6oUqne//Rt
pgNhB5rMah5gu0aMCcfGPslYU6am0R1kYuOK5eOF1Qr/hetShcGW2+ceGDbxdDsdXSHoHdTruYLa
LTCUQxX7Qf+H4Yl2YG6FODqkLfz7Qq0d93Bc/JizDW1a/QWHFV3wIjywkD7UBzs0Rnq1IkM5WY4u
1YpCE0zncgPwdIAK+diw94ere8LfG8aF9SvwOxs7zfAgRBrIJ3EYWd1PE8ZAb1s6xKxKkSYmtFby
x5v3NYu5+MNo1Qe8Ln45OXPTTTYTXn2WHZFnn+RHmXxoeeapwcgtxTynypvA0kmm3qfmuRPDkchN
gXAAqOtm0zCuzSDfaiJkHVzNFITNfJcu9OQvu7tMq2pHJZ9IOqYVdVClbyM/cVjlQrqK7qSK0FtD
TIDdZ0JOj7t7V9Cs/Q+6gp1Y/yPGp7rNWbwjlFVf1CDpSCj4F38eOcnpOHnGCncPBrQqwR0eB0LP
2FcXB7QYgbFdHu7IIVFLFHTcZAVZYS2qEeSJgFqX5fqyS4sWwVAwTuVjODj9LnatSx2bhgty6LKd
ymjYpftW6uoahW4DiTpNyOsvQa0ZCOa45oMrvKnncfmWSJYGyzETCXPSVd4ysqputdcIKpluBqR5
Xzdlakl7Y3vlxgT+SA4Agr3Uu/XQNsL4cpH+Ah52Zq/8lTz4i4CzgE52DdSU+uzrqgnkXAJfMN2g
/RaHwnfry7rqTTyswIytDRM3xCLjuFAwFGLbm/ax0rsAwAcfSRFAYVca7trdrVkEaS5q2AAV6gyv
/TO6gjgaxQupA+I+C3xtcsq9TaZm5wwTfLeVcB9yBVohjt1j9UyGjJXhAD60qsCD5cJDJNv985eq
a69y4qBM//gervGlYVOYXWsV7UaPwFNp+B9gdbI+UsibdzQENRJOJMA32dPQ0QExNLGob9dmv9X/
mw/OGOw77N1rENXc4I4qmr7kRSredrYlfE7RHzl4n1OEucseYwHGiAg2akB3eME61rzoVzieQ1OD
sDi1V5FQUUcac8oSvMQcGJey0w7lQ4i2mYu5BwQaFbLB596/RbEkpsycRTXMVuFxosiOmO3xUU1I
ieoBEcOPU3Xod4hwZUIEpv6AFAB8W/Ex1RJzVEPFOjB78J5U+ArpSEA6l/hT1tdQf+crC0P3sy+I
147Ty+sGdEO2Tvht1LSF+UvToYQH5g7AZjvFotLL3eFhcZi1+Ht9zmhhALTqjYoyOf0Nu8vMOuy7
XtkD9jFzmMJJYab88uQyX2N+Wn9B8UpyAVj+gpu6zr3MlomVpgfyphpn8RNYsny6BFJC1BtVF6Vc
/v2SAdOuqxMeYG8mGTx95wolh/8U8RVDKAIWsd5UDMUXURBQvUrYubx3GaLB1vVG/2qgqXtduDgn
LtPdZ0zrbI3PItF0rl2ynjIjGHMp9F9WDm9ygN9CFeLyWixji7mgFarigsQKZ7mXSPpNzevI5vJ0
pyq7vdV8Tj9tyUn71rkMuf9wr+rAjaZ1Lyx9vChFDZC4kV+JWpcmf8vgVEfRHl94q3HaOrMKSh3v
dvhmCkrx6dyWGwMJ0IyTPxOizsKdi1m9cqlsGz9WGWcs5RgI6hgk/lKAV9amY412mK1c7rEfr5V5
tQdMHQCya/26sSP/T344IKpq6JuRM3q3t4AXWzqklSGS+pw6+Pkl20K+qHa9K1N27Xsj8eM5NmvV
Yk/RZ4L0VlX4F58r6P6mL425Y6IQfrfTS0gyYjcpUgLlgNhAOUTtZ109nXhdKzPO5+dibX/cbqNw
g0VnrekBRcJrk4oRzvlzBwUko2Byp6PPMO3tqHmSgj+DmBm+4c+Vb9Dvgf+GsVLPYBAPXBIxetfH
P+NMMs4mb/ZwbGRpFWKt4ymH7ybRv/e7/1oCsCyRGBfHbPzGV7kFLiCOKyJJ6G6AQ96RdyXCtq2J
4e3k4DI7tCoIitYtqoIvQ6S8ZUO1x/ZIMq6SsKmAV+eKq1obQF6GLNAILaWiwcpckoVpFyl6Ocxg
0lRXj4Jviem6SfvPuij/VKuOT4dDDnl4ehd5TRacnv8U738P7TlU4Xw4mAyN4A1/oEXmo0onqEoD
jzTMXnvhKnxSOHkiCa7z9HSmjDr3Z76MTfmN6OOvJAQ8CJJUoBXuNo43P/KdERHX0XIDCovint8W
bjjSzQnd+LUrTsi6feWAl+fbSI6noqNL/VR70n4nyqXFwFNz44VH4uXaLnMsDIcCQaZkSX2we1gS
hL6B0e1P5hfwYC93dhqgfyQiXg7z9OqcnylRwa38jbH3+NvTO3F/Lg8pcrDkaKyeQW+/YT7Ud0ug
nZUdBsIDQgYQ35Jes8sNfdPlfisiTNxMhKWRzZGRetS/DtJ4M1MEKrzqHbHMkGsp1TZmH5mA76xE
TRV7RkzEzxCuE9ICYZXa6GPohEmNdYiMwi8CuTqMkzfh5EK18KMxQNRykAIK8wzrClKVeThV3Lq7
Sqk6J1kM3tAo9OrkIWqHQF5+tDUir+G3t/9UY/GvAbTZ/caXxbuyrXvyndD48m9XYKiyFCqoyQG+
QsWq8Ous588QJMQ/nHfxkcV3X8yj7o8mAiV6oRmMh7dau8zUV3rAdpblfTie+jzgmYOCSlL3vXAD
R6iD+L8Uv8DLiHF3kElHngCn+7SO6YPXWXZ3mKMMq1PW/+3TaNiIq5Buvk+vaKslwFwktz7dPWKq
6shhDKoOx9hyIv1vW/vYIlOWAZLYd0sNOuadxY0oOFgQ0FXn3/lGlBONEaPXPTOoebFfeEvUtx6K
LRfLXZEKQqWAYbPRz7h/poMwgeLi6q8AAzq1UW0TQN5Fw/dqDKa29+ilbNajmMZj18lqQu9bWtYj
lBvTJO9otEha2W/8W+mNbE62DltB7VBlFQTDVvn5bQ9ffiZNh8rEgM4HrdrpdC4uehrv+bRYXuLT
bRaOBxf8r61hDq/iOSClQS0tCGAuww+C4To6OuNTAwNtq9DrVe5jiR9+Fv95Vx5DwEhcrJS3iz9R
3dgNjBJ2Hb9jpqv/GRXAtCxqEfHRrI2J8sjpiKQSDLG4luh/JAqqOUM2kVf2xD8TlxmzN7Kr2rcL
kWOb07GqBJLpNqBogIPrTsni78Qm16HijzaNbN/7cSTDaj5AEwrDIHNOhRiVDx+md2etJJ7ASZym
pppG4GAYFCVjXZ+gMBBV3bHFmwwTbUUynF1snicHrA6R0oaKDzh0bp9w32Z6m8gfVj4eG64m+jyP
xmSb9fGxVAMOB8f79VH6m9PMshsO389ecJVdJJ5ffhwSMOdc5zRwdjxsNo1qGi2PnQeiwp4T0kRx
j6pgNZf62nBlyafUooe+8/fbMwdwskR6S34UxrR2A7DVEqo9JrYK9KZv4VBKE7dQbcXe3CANauE4
wosGsz1N+W/rSWrkomymgZ3TAQFVLzCaaamDrG2PPRGwQqpTGHzbypWeIDXeFUwHgbz+jnBnQjdy
SbxjFN6esR6x0puXBuX5NzpwxZCEa7VGspSrGmIXt4zVzr63hRaVHMDQeR3Y1vESyUGy7gbvWUj+
9K2eZpoBeB5jbO+0LYTz9ALB/Gykuao105rbz+/DPCyv4aca0jpSU3bCeKHEbmso3zPdNsZE4wO5
Vgs45dZUL+O+05yDmbKohLEwXf4i4/btBODlAXzbnKpqVNGln7cluKc1eYahUlVkuIwpTO7H7m0F
dMMCRSHQ/b50XjmgDnxuG97+cXQ0GrVZLPKIhc6o+Pu4eMhAYgkrNyMYXyfL47qivkB7VX4CMzcb
JgFG43K55Cc2CStCozSPeqclGI2I/BVCLxinwr+uSnGVqlr1mbvKBs2UgtXC0QjkiTwwuj0hvpBY
mJHkWcszLaEiUBcfBHpZ3tdz+c9FxamohmB4gMA+hSZ/jM93mWwUpiCPolXZouiQ/Ga6OyWw2Bea
FTYpIuvbLl1vw/UB4LfsjO5DZ3rtbazP+8hYsfEjRTYGzdmOFZk3hfl1ZEfITn4ibpGQaKqklSt3
DGZipzt1TE4AWBTnv6ZI6pCwL/KUCdX2AWFzbGDjetIAy744Fnljj5AYEdzRiCCZio5AlpgHb2fW
rcrwLWPzaCEslh9tUJZ1PB1Irr1OROzAPw/tpV4jb7v1ICSwe5pk04nmHe+HLTz2OdjquLNEujSc
VCjtvv4wdVTVqRLmGULvnQy28CtoNaFuZ7hYXe+XtkR6a60hEAYfj/sCMc2ADzm3/dx6IHFvgmKx
njikqUVBz1mNJcYDCHHG2K4LChbM7CIethKMmAIyQo93jjhUCjU4bEX6F5thG8eQxJCPHFG42b1O
lk0UaxSzzouEKjY46QfDjxWymZt7b01sgjX0HIV1MZFLLZD9VKkhSK6wavHasUZvIR/q5HUGaEHo
PoSp+7kEOSwqJC6DkApLy5W29G8isBZbb4aDAfxdQHsaGHOo4mymzB7zzvTBj1PAWsn4GfdMD0HQ
c6LIEFwaM2tRXaNE/tc3D1ha4/6mAhnHy3HQD7m+i1OhhfApJhF54XZ30Gt5OZjKbx3SJ9WkD7+7
Rc+yIcc/meTADwHYZXOjU2Zr2T6h3dDoeOR0yQ7pvP2yt0T7IKRfh22u76oCEN06r4+2CgISQKWV
S4QBaXOa1trnWQDSzJf3KI20LCrjxwgkNLzgtK7gisJEMTsBQtHsuPQ5JF+O//Q5XJ9JOOqAgkIp
UYQ9PIpeLoJJv0UUwE5PATVu3qnrRPMoSWMJYo14S57aBpg30tDeMCwkfOtRZS5mHVanfa4SoXib
AK0qBFzHxSt3XAnMHNQ1R77O4TsZxN4KNbh5gADFEe7XSMmRtdk9nt2M0hcYCTFxAqjj/JB9/5zM
l9TMdYkaNL+QmoO6bobDeapstGTfDkw028j9yJxXzTW15OCNnoZXjGLFfth28pcz51oYXqQ4V4NE
3/oDSG/O+uuLP28a/UinRMh4J+TQbv/+cB3hTsZuzOcDoGy0omnvuRVG4j8IEhdOSu6qFFARZ0AI
PjUGJhFSGOe6uAA+J/TyHDklGkUcE2IRInU1gPdMf/izZyuIZ7fS5sVijEG/bTI6WTVLdkNB/Jsc
b7WQUwQgFgY97xq16vV++B2tKUiSBIF2v7ymZN0zcaVpqR7hA5NhTqU9530fN9rSEjGbBXdr5CaM
qumyEYPwKYC+Fc3Rxoir9x3zRond3VCjM/biXxNL7E9EWjZUUud9N8CnQi2H9f+5S6pJNRUoHOVX
vaofwxNhL9OBhOO1SRZ+rAzTnFFo4UuIN577+4KkTFTMBQw07Iv47WYrrAb2Qa/NnR6tpoSRNi/+
4675kMMk4u7x+1RfOJsWOT4OePk17UBBfyoH7XV9kutwccQd+3PKMavMKY6SEHq4wqe6P3u5Ghx0
sAqewDUVG8Upge7gUHfUf64D6mvPU9aFu5qfmBPUBfMScKSPkaSB8QysS7Z3X0uAlUe8hTK8Tdeq
C0IUzkEjXTS4wO5ipVcopTt8PD7S1vZiEtktu2iOgxrwP+EctgxJN1aztrtCLN3rTWWOZfjGzBlX
aQ7XP6TFWYmtbnUp4qeyS6hyyQaYneXvE1GLYuhJGP8iVkyUqq+ykLpdYpZz0jDWjPkavIkE45e1
Kk2LSLKrK1ts3eIXX7Dn1fmTap5m1dxXMaeZnsVQf7Joq28GlI4JkdMN7Q+uyAF1kMVt7Yj3d/iU
eu6PFYTYU6ODJMda5d2aRIlBpONDX67GrPhaiqrIqL0blpWbpbovEuNDcrtc7x7jQd092orU17Jq
oOKkfqgqAOwZJPwCXF4Gk8opJHIyVbYSnB3zPz5ZHPseImIjSEz1Ig85b3YY5dt8Y2m76H/rvEuA
MApluoEcknnwVzInnU7WUPdzAHq9sKzunW6Zvyrqgo/0FDV8NYAwOhffvZ7iYWp+TSDlXFTjN65e
VzGAnTEMspysZ+/TAzfpMrI4eYuamGWHe3+LxcNaPLPHGoDdARzBeFMq9NL1F8yxmd2tqRMfpArm
ZG5rDRsgfUEcSsn4Nf47OWfN8IPOSa6qIZdsNToc5ftvKVfajxFRwmewgQMPdAcHekwT04czmG6X
gLAThkLIEtEzpuaeSvIooT4NUzXlbHN+OuXYMuUwJ242kOKB4mF5EMPb4P6DTJEGpXhr145D+kSD
ylptsxpbQRL56BEiz7XYPFHdKWUluCdZ1tMwSoxd0aPBonxHf1yhN3WTcDx1K5nLBjwIoT6aEYEZ
u6XfomjvkaW3tIGVmYhQn5HeMgTn8AzRLXoMwI9XVTs67Xe/6Vj6jMQzh1T4J86LolsMmq3MFWxv
rDLN3PrBK1i4uTpAysnksvsgNTX6Cqjr7FcgBikYyYc7HiNDrZN4/q2F+CVwFlkGflbfXT+JYraU
30otub4CuEZ4FQRDt2mOpTGwHnmz883U9ntmP7yfH1/Rn35JjBN82lQEQiGRhI+AcZYbXCSecmkg
eFc5c8gc4ZiSPGpUb7+Sm+Lfpz+hTGLAAKvM8YZ3rdCN97ErWhIwHxBpNkV8H7zZBMGoPebA6zyF
IORe2G5lELpGnpTc5LTZWZGk431SgTreyDOW3V3bWK9zkyg+LuqylkVDageFjv33FcUNgcXpv70Z
yOdqOo99kqmOurolI/gSZO9QnXGxGbk5rtKkTqTcLKfL9NyKD5ZFMbav51/Fy6kiY6cbcTATI5ug
Bocf/jq7rf6s37wb8tLmzfxVUDKwHiH6B3tJI06uCzS0V+aUKq6v+gXkCHabfdsNtV+1JqCtEzJX
QF0F4Coe1tZeN0uYEchb56y7fO6rOtrTEeLWXlrHHvYJvE1CHKE9FXkpAK3bnj0NZ9bo7l+3f7XL
byUxDL67sDMBpG/Xge+yE7hydPnIgYC+iV9iW6EiFUheOqobvQElaUbypAPsqcfC3HXhxjNY+XzR
P/V5EfzN9tqzWFyQXW238YOr+1Ej0HfEcvyFzj8bSCGl+H47j260Xp2ILOvwg1nRj4GsJz8tLuZv
m9hYCmq2KdVC12YbjGpJ9AH+802UnxUk0Tqh7P+Gw+wRdduhCbs1K33v/nzEmgU9zIkuWZGjByMG
BZAWHzq7OshPYIzegn4QPnGeWBA+WO4txR/zDz93Rsx96IwFWCXpG3cGDrR7E5QzCEQW088nHFZA
mmzoVliIIJpZqUswagXDQRyveFSSwqjmBxHQ2sblYMGGXE4FOO9bQSGLuB0xZowAMLr2cwOAphNz
Y1iDLuoJjAsieMDfdNSNQnrIAx3F4zeB3BmgKN/U9tFkQxgyLMvAML8orB+7xuWGeDME5x+zQiok
1SE6uACIs68SiXZ5mc6bgI/B5sdZxtB/A+boDEBRs4zoTSfeVvPe1n1blPHgEtesUDNEzfYU5ry3
scBMMyMSK01rJex3SJrHu3mqBbQw8ZbH3Z33L3Rde+9nbsU+bsS9/r2L3rcG3D9/kfA7Av6w/6YQ
BpXFAwNHD8igoJjvHrA9YQQ37zstxc2HtnwseV/zmS/Fp1r0uGkJ5f35ZmrTLmo8Rego491qigJZ
46fTyRiecG83NXHBpCplImeDhnDkSoE1n21kiXqYAQQOE7tPUNwjg2fdeVoT0/jXH/nRkLRd0ls/
6t4VNy6e1I8Wu55bAcW8oOk7I81Wz1vbnpQevjiCdo/LAst3FslEx560odXFfkGnK1octFRctI9r
xta4a9Z1dh+W3lO3iOETjzWBfLKDo9tuuHYaLav2c61zXB+btB42QwuX1Kr4Sc/kk/9AZUQPq+CH
GSm5+5JUnayf76dYcDFTKUFX0aRTb83ZAuHW2Zbu608SY5RkDOJy/Atg39OqAL9fJwsujvczkN3e
lM5eUsLdwmS/d9EbauPWJYIn136KptJvV2nSQlTbnacTQuLV/B4D3uImd9itTa8O5t4VR8M8chc+
xGyBlvl/McXV0LjentLOGFyXSvTFcpnGJ7E7QiEtUN3yqP5A2p6d4pwNYdruW30nSRflM9FQ0/c1
4emQ+2u+C7DgcjZe58xOvvrrI1fCU5zxgoKPEFnVcBi3FjfG01v5erKIAhCuXzI34dHAY+Cva2qq
asrN7qRxl+ClcXw8R6MYWN6n50CATKGqOOiPa06NMrN2MEPYdxdxhXijjdK63oUh3dyv5zmNTLpk
qOQH5vRcPRGHcHLgsXbKkaSNFMW6UpiWuMVM4BLp+3xh7cP6Iyvc/Iki3MrQi737xd8506xcTe5y
4cTEZZcp7xT1tEnD2lKSuZ5tVVqzfBQsL7GXM5cKQM+3NUjteVjdJLGwUDtvJnIhlDfzlL+dRYKW
tX+sTsGL2UpK+rBVQK7B7Ov5z1y/+YnSGqWxT6/cA16WZxPLYxykTY1/7h0ZPT6fCboUs/M5rGI6
2gxlYMgR+1N27Rb2wq8pLSlgE9j05G67l51rdbEUU6b5uQQQRylMSQJgXDbR4gEBLLyT9Y+Y0NvO
AJ+GOHbYYSXx1Gln0sLAJylhpRKaxNnMuMXPmi6fT+n3b9k2zEkVM5jfQOonUvODoQXNLiJumwtN
RuR8Qe+uEkJRPoTSH40MFzVEPuTTBtpcIhSsVakqv2B5xMTdE+ViA3GKcETFfviMOywhiFsWRMJG
ZHW3w98hVB0vDH85aWhk8460AkBKpsm1dE8M8im0IcopyF4AlWyR/PsOyLRTW3U8bbIpBq0xwV2/
u5+o5WAWB5WSmXw2RktIn1CVRkSWXEFhIzf/zt8bLKnZwpcXg6nlv5idbmZabbf+tvkvJFhFMyxk
xNzzjyKIwsFW/joCEv0/7Z7CX2yIbo4dOEc1DWhdFGss3GVF45fumwQnHJC3tXH+2nqDUzMgV1MZ
WkbGehu5H/WmW87wXoCUCXXXZBcZvNDyIITAzzNUXQ5g/7E5GM+378LlwM1tiyXdjEg5PixrBmWa
Ucy9H1MG+34u65CE0aE929jd9prd7AYtNnepUAZE136BdX3QFLF5Nj59wEU4kRql/zj4X3lr+PpM
Q7LJIBhbJoaU5Z/mSOvy+LWtGwBSFrUgs/XLgyEZmUun+cslGoFxtjyg6W9F8mDZjppm4ANgnywq
hoJwOsezJ6BOrKGOjWuaQ2e/YlIBUH0W9j4dkqXhdLekzWrFfw7cSNKgOdt7/IWOkB68dWLvqz/U
KPPXGsenlM5GsPCM/E/wDKtKQFFdPBE0v1a+7D0HEGlIIky/Fixd5PrwUOBsgsw5hbgybTLkJH8y
dwmAtYXqwCbmTXMpwzAK1HoWWJRyjv7UDghJUK4yyEWambT4VKkvXuS8MCLkXT9ZYnoJ29BmEp/F
DEb8iLte/E18MYR2Gx4KDmqZIoc0jFOPnJp5cdln9ktPGXnfQf0zbMHcis/SujDvM1Y9F4rI5dyx
qp/Oj47wL8dbfMn0HQH7Uw+YWiagsLKpJzRSCrVWO0TTTuId9BdJ3Ngoz8ZLlZMFV7NEXqdeu26i
eLNoqX48re516FvS8MGpTIvvsJidMdmExVRtVQt2EaplYCBQ6pEs3+z+a+wwUaGUC+Ib0uWte6Sm
+MNifz4+fgdy7KO8IZ/HMmobozlp3rkSlnzfh+B+WdH2xJ3v8il4hOrcylTn14z6IgLnDLCXz9w6
JjYxshMYL80nExrPeL19ojih60rbn8/p86+m1uiGjnTdwVVbvCa1bXSSiq0BRUM+9E1MNPMqL294
/t1mwrclFSZEqyp+91vyx9IUFFrtRI86i0/kQS2yLhCfgOFlvXTVzCWhPorDlKLuztq5r4MthQdl
dxpOND5JBZL9ij9pgaquHwNNggz8eDboWxPxDjx34HNJUw8G+EpEUNTEi9k1HeuUzOM3+Y6tsPgB
IxOwlfjhMj2TEh+1kqtCoIRW64HL/UO6nEuyPEbLL5A3ZnJF1aA43SoYuk72ys0btWqWnD8AEnJs
n7mGYWd1/sACDZvgPNwh4s8vqUk5BlW28US+H2FbtqxmwefXR+jNU7rmhnkLQHpXe9tR6IQrutS0
Xx33ZQapdAG2vjLlQQTU99u5TFGXlvNnArFXgnOjcg+Pr1YAWSrTo0RvPxWkR2IEIRdqXbd1u6fL
+I1ByyMHSh2KXNGAkkcCGg9kSnnyaxFOGVvdpwtSC/4+ESDokwGgFM+BglIRNCS253Edn86UMJBB
uURhLWmfhIKJcXvD9Q9iAg5aSAuGtTTm8xV7fEa8yzSZJZ09O7Wj+S1/G2FKqBy0vb2BREK4Ygbe
/Pn6ohzZ78EXRmh4bs4BrKQJwu1gDpADOAM1kp+2hlpeo0L5yQM07OANtUhzE4M9q82JPJj0NgC0
8rh34CL//N8E08Kos1O4URnqGTDrycAtJzUqw9/WW967/9Lef4pVVp4lfbW3nsm1HQlgko5jojMy
J3RJazDsJ4XfK7ECOigaDVcCLQ3Lpt9TYFemjDy7+g1YwY6cFiVs9cLRTO+cnO1fG5emO7btlGDW
626EeucIB6MylnPu+FmQasN1mNXIRJYLqiqn4im4N+lkBxZ4M4H5Rf7ZYxtv6cH1NLGxSN4i08qI
qhXXfd/4KHNT7Yo/WEo7lME1H4EKg7cH24FEkwOvnCva9OCEIQ74cIgbaT6xMeZM6ipMZBBGXM35
E+uZfdm95ruTd5P6yMD0yh7qFYws4Z9c1K5xYQ5ZKgFTO3JKxFhgwLMKuzxCpNQbZYOjVNuXmUQs
ogd45NhxUDriGSJZ6a5UbKPWyfJJBtCyOrOHh+YS+CaPr+Osomgz1UPEeCZ4rpmp1jgL4xRqFgaT
dwo5l34jAW0iN4N1P444neFRZiRGh9hoB9LpRYHF3zoQ8h81CstJs3aNtrCb4n40rWJVKKcpIsda
2QPrz2xtc8Hg8YrcM2PeL1PXratqjH70JK+Nz/YBuGkYTB/8WZIKAFxYhV61pxV37khNJWZMNzEn
+oxALANnCXtNvSGsIaFlDIj5g2f9+pXP4ME0/QUHKOLaBpMgSbK2vHRLq93w0XOZLmfShw9EF0j4
1w7cA6NsPiCea8K3DMlCZZjVme0LrIsOp34VPSBgv+5pW6e3CkjQWJu5xK+6Qqh+uU1CPfOuZ8U/
HBNaNmoj/7J8/HdY6OSem9l4xQvdXROxnsMQsOn4WnHX71gRRa9Bt9hhzU+90fRtuH2ime/KjhQc
hEkYuDiYZCMPCUtNGrqtlbDQGctXigXvxczUImbMAHhXawWE3VL5fMhChOO5N0y/na4acXfEwJIE
cz4EymZH8U9uhZUoylhs0N3ONDrYDyMdWAuC9aGEY9d7Bz49xsOR7Bzf6/Mo13nCcOgElt3LR9SN
eCibkWo/8BoiNR9CXeXBXxMVhJ/2lsXznAKsn7Og2m892JOUSqezAYUi97K4FkTwasiWk1TlhNtk
CUWUUh9LFyDDGTExMLS4LFzrVKsNIvKkxgoAY2QIubMhICH8ib2AhzGzkFWcpUROa9misxKtmYs9
TJKLzMDuBm+CaYWmV+VSG6XOWuOavPFaC61afKNbWz0ANV0W8PpF3PQZCGTPY5UA1qbwVCoRO23z
ZtVmoKC3NJQS/THvndUY2KxWdzKg/47+kUZfP9oUluTabCRuV+9kh3jtOh6ehqSa/RcuG6MrVj0Q
reB5RvdZ8UBeW0MA9+JeRmR6zM9ZSjCWjG2wc+8L0ZK6KEzsO79Pmp1o9B4ZH+zGIru56RHtgZbP
+JPd46ueKewkpIyjiQnla34Mf31BOPW73fkEQO9BqzeBsHYeuYimhWC8ksCmjunJjqaAcrYy+ovo
dGtkoHJzw4VjCJffO5u0pSlui0rkZcR2MDl9Z6/VUdMacgZqTfK0uwkC182GO5kp0vHMrRxSnz5e
LDibfS7vhALj+8H7svV1XfW5Tz2EZOyqLjg+aw3SM/0h1AFukyEbZfQBUCq36xzmzL2xAGExeVhI
jpLJD0u4lr5Tuj/MCRgDXYMSKZduyFIMdvw1eSGSQcj0ruTshPILR5eh9Dpxsp8GS/5YmMl0v7Z3
cLl5ebHxKCQUmiVF4aaviIIwFHe5uZt1fjmrwvAQCyVfwUwQRsVdlf5CfL8wT1ST+V+tAtCfL68t
sFKDHbg2ZvsC4hUvIEmtOj24nH1DOHDf0g5YIFdYg98x1FuC9xHidsrq6k3pz7FLLgQ1kXuzfg9c
1RdCT3GQ/19Vo4s7oAYgktJHPpLDmnfTU3M+V7PI18ZnrozT6k9O3TSMMW2+3jYNrBBa4S6KY6VH
jhA0UrJg8NnXq3XY5gzYZFcHfhydslareEaWm7GNkNUexB13G9w3eq3hP5Jo8yDjYeoA1Ldwl32W
cbF8JzaU5xsbVxIp8/7e9Xd6WYHUHdyQ0ZzSbVAqBlgkyWWBSPEUCrrzq1DgszBLL3/GEIq65QAT
Jl/h4qnlWW2X2ID5DLNRkkaV18mBru+ry5pId+lKMBBAff0ulkuFcbtyke8XiMS7hAXy+k2qflu8
Gv8419BlEiuKfdAQ8dUTGF5AfCLfXw+aotrvciofBmxQ1ibiCDaZqHkFWY/dhWDK1tHxhKUyj130
gNNk6O22upA8l9m1mlIcs+dtxfkLGqa80h7YQ9OiGejUeoonVs1Udxv860DYiPnzslaoejzBcCuz
SkEGGeRNCdbwEN6qrbHzsDe90vlOtOkz2b4KXZtraY7/AgYfTXHxbKn9dViJaChv//cw4/eXEgJw
5y7Fd41t2g0QRj8D2brCO5K4OKGwfN24IOXWHfQAHq4EXVm1enNHn9rnO9i0GslaJSAHudU9iU+D
ydQ30U+ZJN0j8kai79I82/CIAcOR1OVn24b9ZQrP8PT5WQQRRI2cg01pm9/kIwSysQxif5hC20e8
w7NSYWXvg08FRNaL1W+aAqhPHL4mIbmj2Oe42qBg8sNCe6cT2Y7X2E/Lf80cFezJ6jSAsMEJb5Fc
qLqbgeP2tXFfQCwZ68689GfEhOKi3sAUHFhtifpNneJH/EAQaMDqKXUKTrLv2OvJ1TTyDXs6Lmic
emoXCjloAPOvezuS1W6TRw4l4+SZnfCXJtCnxaVnhmO4ZGIG3ZGbN8FnD8jKHdLwuUM7Ct7bZPxZ
SFWD+WRpEbCV3jtS7leRX3Ok/47iA7redDb4CfbY1vH6vbFS9tZrR21wmi1qd+KWDhJiSLLGAw1i
Ts0MDvlUTpKYMZJAXcz5wJQpEJ2AE58t4sqGk4NEI40OfMR6v9ouNI4BHF/uvjmlhP56jkh+p0S5
k37sLBxadeqc0uCYSprE0orHg0deoGMhfE+BT4ysDBQAl1EaiYNahSeeJgkGkbE6yO4K2OnO64A3
iKO6irnI13Rmv2UYVTHXXRL2gUj58UuMAwlSISEASf58PwqH6LnlSX15Rpylijxx4NM1AIkgUOe0
Rdlc0gG/OL9RjP38O5JPldT+TN8W3XyzkLWSl6J6ufcwpM66um57dXBuYUdaHZpCAzUN+53cRhpv
eEBK5lZywXab0IhF9MKvCk5c3VNIbghYVryLevR1UO0l27RraTn8ZK8vWr22o5qQZSC1axqySBEX
78fVVllfVypGxMNSBzastdPUTR0e3RCCd44EZhjsiLDNUc+HPdF4F6KNkMgC9IYzyX+SM62trm1C
tA4Z7yGbEJWueI5wkvEg0FnLc/4dZUbnR4EfVkR0MBol/gVUUtu4QA3py84/T79VQIzfvHtsbHSR
2knlxjQ/tPWQOq4DGU0jd96Q06H3X0sxThnFA3bjWJ3ZyqOYEXjgsMj46jGisuZtCKIPMd2MWBRW
/ZozWMXyOLu7OSWgDniUA1/qnf3DHj6DX278w04OWkwZYVrQ6kn3eAu3ZW+Gls+4pgFxFNZleMvJ
sJ62Jo73YF6izkQpmqKfPdUELOcG2QIVReQjX/oHBbI0Mj6hHTsWwG/axK2NYYUxSkQCxjVn+VFw
zJoPyQeAheLOIOjOMavm/TvQFPLRVMNr0X5bKlb+MTw3xeXUFtW51O2f09GFitDbzT/cideNkBgl
uXuKKYHk/3iX/XkkSWaii7vbON6vNkjfAMnJjFpFEaLqPxTx8zeSbLp9EDeenHgvrNiDs6p9CU+m
excuMKfPpYgpgcAW/oYd+Vsm+DoaVaJI5KwL2rb8L5pOgzMLrdli8HbAnjyzFuK4QhaXk3lpV9ew
myRr9UHtkrIPVmfH3tCvI4tXQ0wmMILQzYi0G8PpiIeuWd76c7oJ/cyAGKak0u28Yn2ENZZNy1g9
uG+es/xBIhPFaH6gGqd3g1RenvT5TM4bV1z9Fr9LkY9KyHNrNAAnEqu0vouli1+M3jZHLnYoBTg+
ajq8uCE1TqNZVSO25b5NrEYHrkrqDdeQbGYfZ50UjSoJess7f++TNT33YiGy0er864M92b07tycn
FM78rD5t5hUz+SA0ftJSDkU8gsgllsJ32AfwGdE4GqR54ryCn7WnPj7Vd7o0Ix97iWDZDHmraMzn
l8C+DsZ4tH93Of1he+0pkcttgQ1zfvISneAXP9igxiydnaTopTg9V0zUi2pXfnhA4y1/1MOy/TR/
QRqWI+2/1BZ56KXtGSYiHrbfM2ql0Uy/s/tuydSxw4pPKKOiTHGGdTcDvTqk1WdRjLRps+9QTSsd
LuDWIvamY0J00hf1V4t2ag3R/Vrq4HHx6SwtJIYi4qurfeQ8mz/7ZvBG5+X7BEjGiUxPlhuUhVgL
K4HPBBhI08OXzemIeQiVpSxorescMVKjKxF2EGa6S7Clg4M54REm8I6QErR/xfnRAf7mGq6uISCU
jznP+7+EHQcke2eIrkRc/UNCxXTy9Lw0K2MJThCwx+LhHRxb+Q1B2Y2GitoySukAke7Ag8Zf257F
IB+l8D938B5nB6hsdQdcS266XmyoYe0x6FPHePQmPUDsQy1UV7Abi8ueQe0FEbsYv+kuBQ2aPGCk
tRlggAkuuTuupim/QCE96V2ER6qmd1cHFsqI3TAI+/rnH1icK9TJLuVx53V3+D+xX0ql4SaTFvkq
Yup5w0IDUbNzjK87g3V8AHqUI2XAHU89yYqxGgFmTe717iOLVk/6++4YIz6m7Z2PeWNXiGqRTXNn
zhWZVnyqjsnS07xUcFTNoe27DLQH6xwlDMMUAK2AX2iKfq4g7INcNGYGl8Nd+PXVQ1wPYkc5bmYa
EEAw2gi+/a2vSP45CRrIs1a4TyX3bq2DP3nAoUJ7yUq11D1mJWdjrniF7Tx0IlmHgDDnOVaxDOPq
THjrfJLfzVAqFzLw+Cby5/23SVlVE3yrCZTTXWMDuxEVQ0dMO30sMkIrB/9tgXNWOwPDdz5LV2zl
+mepiuXorFrWIcJOJILEVKAh/At/rC5WIIW+IorIbvr1lq3vZJ8K0JO6zz/bQnoodn3vtUuzjwAs
nzXrS+RsLiNxMhAbVsZRouQ7Eqgbq+HY9yY5+BcfFV/nRPFpm8MQUzsuK2wtIgU3wQa2tzduaHiw
bM+YXmDsW2MB72srjTwGS3AASgYBLQr1FdSvEPAFN3hd/gsxbknA/Hm8xx/w1/2EySaOSYpCJj25
jPvzZhWVkiSuO9PoVCLw0VejqDhMF4TwF7q6QD/4MuicdL1/RppDKgpuC3t/DLOPOyg9DAf2UQH4
uCNNLevVFgxdKW+UU3kOaH/5ugn/SqYIwdEDt9YTFf2GlkG0OG9+XlEHADNkG06N5aQSvtzTW3IV
Ygy35qNuQN2fQGbFq+czDMt2QjO8+Rfq3vNAoyPsIYYL+MXimxpTTXFq8B3Yo8XyJlkpYGehT2Dn
2fBw7NVlkNz2AuCLxpFPplCHq4ipsRoxBCyvJYcwYyhYT5Jz6snm+l1hMmt3gkDSWrBNaqSJmQVm
d7jkTpK1mE3iHl4aGdlac330EtA3JJ0pR2E6yjcJAQmN+R3EsMpVTpzCh0CAlkNlS18bh2SZsI2v
69KdAk/S9bNrOqAS5YDM6T+O/abTpWpH4u63xzPJeYrK/5ODhlBFDljScQ5c9efZISEKaFeGIWCq
sMl5J9RW3ZDKFOyC3iqXpGnmMiHHq59L4nH4Mi7Z9Cw5D4850hr/31ZwwhQTbSrvFy9BPcqlLWKc
O+0PWw49/vKtNNcljswQElSOfesatck35XGIVTZj8yreW6JS7V3SdZgw6noJN6IPQd5lwz+h7xtU
mePgzYTOMw6c46AO7IH4eDCqFUp30mIb8HRb1wqMoBywauxa7mh0NiiY0W9+mYI/YNjvwpPta9fi
B1lRPBKIpLHzucDfbf6fzSusXsZamBOHGWBJR2bqPYV/UxZanSJqh61E8hq1ZEmEzP88IU+YKwek
R4sYD/yhJ2r5JaTmadYIEJcY3EhntPchUGcNK7NhVqAd+70ig8M9GMyrS1kDcXvdw7RvPjMQt3zY
uPQhLBGb8KvnpetffdT+NCpDutfh/r2ORdzeGl7JV95ogMtSTvTPMBYJKPQAPTOxutrOOLwakt+7
hjbK2+jV4Chc0tECVmxcJlC11sfDc6BaHbUDm7r2tKO89OrX/dUQMdAeJY8dRZydU+y66p0APlsq
a8dcuGmktWbg2mfE8SCTmYTIQ72m/zvIf9Evn6XrXNc1+4hmF4ysgcGvk9MU4ncr3K5J3hQJK+nJ
UptDHRU8fb4Iom9BtiMZWPBUjauWnCa8gkv47Z2DQGV1mk1WpLl+dMNsGHRt4bf4yYmKbabbm+bk
INaWDUKwnavalQqhv6/XySbQAvGzUzqHfD/EgewxafJ7zX9/SI5b6YSfjnQe9XJZpzYVtOFv7jQN
A57RL8Je72vLvR5p2AgMlnV69CTgqHJ5H3xPpuJMGAFtt+l/POtTkvTI0lrHH0Vv50F/Nz3gHdop
7ZneyCC26KFSgtGZnGADKtuUj2XGEqouHxqntHuyYgewmwoZcL1NgaKjHxaMppqSW4G5+7ZjlogJ
QyS4gynVc/uqlwd3w9xSLwwdMoLs4HtRDP9nOds/gpxYQmZCyTvXLiaiJpDZZZfF7pF+kR6TWwOo
D8pZp9eCtNNJyhE/LYOw1qXDZnrAFL7bcy1u8nsbJHCuIoGOOgcIspa5H4eiP8L+rZ/OKmyNE/um
fOK3jInE2tAfN7l51pbaNqVco5OarfK9LBP4JDVH6qXwHypnGzWUTF4nd+nR6PSkBKHDwL5v5Rg3
D1d5ShRm1GRRrLzEqUiq++xV9MRR04ob3DYXsrgfl95C+FUKilOJxbJ0YWy2JqfsTFsqh38xg+Cz
N15UrllrCKW6ZBGQ9aFKx1MD+GlcV1m7U/YUVGgzgYjoICFpiSIWZk3zEZ9oyQKisoJuuYnXwByo
Dk2/C1wVUq71fpCrXBDhZfRewz6I8ltQ2AQSvHnS5Vi25VRERBXgm5bmH4o5wHMc90A1v3aoOac+
eBicZeTEVV0yhPnilYAV6WrEFoaFb2gf1Pnfv9PBq4vjolyAfMXHW2kBlsTWtgHYrSBMlOn5bLdx
S/aJbf0IwI0dgh0UGCvjIbxdwtTBEweQazjOIhM2QvfOc32ILW7x0XypqkUsdIq7WdfG1y3pBwmB
Bz4cGMna7MEHprgVw8iSceiIRKCsIZbRW2Njv27/lSeI3jmsVzAmeg86Y48nsYiCgkkDkEGq3CKI
MpGyz6G4qUW85A8JCLC2VkRUfRHfUd2VB+p89tpvAtAkTduBJdBSoBpY9QJ4OPAB1qZHi2ay7gAD
tsvrsKuxzjktqs66vv0cVwybFyns2/Na9J6+slpN7z1xjb1zuL2BHD60SVdKitt9TIE4pMP72aGA
3fGpG07gxgRTOkB9nkjx8J/4AI1ga6LSmbSwwYUKvjnmxYfynwroLQps5ZcpB5+iaW/OjOWO092S
F90UCl2yJxBpf6oJYP86Z6gejxn73FXHrGHBcQcYvFrwGv9AomkIR5HfoTO/ymK9DxOfqhVpDkdd
LUQO2OvNKjW0kYGkibPBSxK/UbDyA6ZHL1hBQyFNJsuksCMtzF6Gd6to67dgTwk8uFK5grAJnC0B
xbA+ss9lzaIpjRPuZ+nqgK7ZSk7ylHIcHDV4eX3zI9o2oCVAavnY8k7nPg8pQJBB7UyKgGghiRVW
s+UlxbDWGAqbtvAk1z8AdMBZp6F2uvjFiZezBbIxmtOdKxFGOMyuOJgHTeNfLkSah6xtwnbEToUJ
TB9ErYQJwOU6h3t7G/SXKCTB3HZPEedzB7j0sGakzijK9RJTHvTDEiRB55BymrgnNeVJlFzsLE/R
nx2CWvE1bvJVs8Ql4BZh/EeuvaBz5JnoEX35Q9LEmsUlioYYiv4XgsKjOm9N9G4CYL8jjzH8/dPD
x7VnEFOsvwZdqPK7vkiJ6o+sSWywpEMCuhJPI8VpTl/XqUxJ84OS8bod54Q9olB3uTKIVyFlKaPD
O2bJZyhPYkZqZ94kY5y77KvhDj6LBvu/DKNnsYhTwmJ16PQOlimKnwwBB892lQXgeTNqTKGEZnHk
Pf2eMFKfA53uiJYlb0xTfjv0OBA0qUVaaa+A1Obv92CQOwA841XqKxNAJJD23y83sGHfOJ/FmEFt
Se/b3hiGqTaVfgOyao+hbLWeqsN8az+GLJfBUzLOLO005TPVVr6gM9Az8x2DSfM2fIAB5m/gwR4i
UBilcEpud9zx/gckDqwjE/DD3f8Njw/DjixCEdi4PbnA2HqajG7BdyJzDDM3xmzw/cOOU4Z2TO/B
+SfHXC0yLzeq1utaGu0DFUVzahfAKkwj/geuniLtJb082tF6C7b2V1OMGndMPpzDDsccBv6Tv2v5
2WcymWLx2YbJwpqpzuhpkQvnQ2cfA49OJSnQ4R397F2Xif/DBz2JZdZ0QSYi+aPt2AkCEdCDTeK1
W5D3yPCY/3WBM2IoeJzR55aIqg64XPtA9lzuawlGAxAb8bml6Z5RFshD06cd+Tu0e3oTiP2AkJNY
6KsEuCBvyY0Eyvsra8Z4rBA8ZabBIHDRxcEqM6BxupBhlRDZ+8ATP3I2p1iXcOcDNQ2IBIDpmUcz
RmEowSLO9KYwUqIEbSehNF/4cLDHQAEa7FLxFwYXqS/jBuZBvFlpga689byuAI6ZRiYFJG0fZZb4
58Un1Y8tzyDk4Bx8VEK1DSWrvJGyYsNmiG+cKPe7Mh5gYTXFlnL+1S8lpI0ueii0soHyWpDxINF4
gcVxczhEnnUcQAS/M6H5fDMocQsqTftNKUJ5hyh94GNbPaJS7H+eUS9kNCECDt4CEybrh0jhNWoc
aTrZheFlWKZewIAWgZ9G9Q2Dj5WznhqAwwKf8E/8uafq815wTiZ63O2QlILOf7/A55eitXvnau6x
XzGGoZe8YKD713TkEQ7Gm/TcBCBHG7bD5aiIiIFVmN75kDsnVgH4boRoJexBx++BAEZcp53YlEN9
t3OyceU0tS00sZ8nLrO8+iPtTHQWSMWXP26soNniSbCkoUH7S6IeYhSzSv4q35FyfPC3jcQWQLk/
WUDdGbF0muZ1JSgIdAtQHeRm57VQFCrvUZ2wdWTuQEt+4ZNG3NMiVVPrjEKQBsNhQmr9tKO67NPR
Ny88XMSNzF9aCmjuFL01F653LaUhbvWSjX73J4JaiCZF96ycjG5kI7ZJ3RwTSop+4OupvM5GZywJ
YQYO1XicGXsgFSAH+4SSa15gzNCMQ1mGypK9Msk9oo23szjQDjww8Af2wGvHaEZq3zZG/JjPWRrn
IkYakAFNiEbyvC6bxrNlVGuuWyEqzo7pk/OcyY0x/d7tda9kMDz9mIOJ2kUBs7sN0UrKiO+owliU
cMz+9J1zGKB8zYh22S9AwQzShlXmJpMdrH6y+uvNShxI/gw7GRIvxRvLWxg7PJjGvYeacQrj7Qme
CXL7dQf1lJFx3wpMM2xLCNhGqSaP7iXIA34smdMvq9r6b+QN1PJ3sFT8YpSgU9mB6Dlrnl9ogL9X
3fnTqUehjrLFTdYgezq/+OQsmnGJKF3JEtPexEJwSQnq0k0q/O3YFxW+xaUyBOV7Wb/+hn2xlz6k
VESL5W8IgVFWX35K/UNX+pmAQJ0DiCR6IQXo4dfHQ56rTBgm+IKnsEFK//KjFqIDuyZ+0W5s6e63
728lXuQUTXQHsFXReM5+GuYz2wniMNd1rX3kpoYN6SmEkKD86+Cf0/rGHBh+KIhN+VoDBbVUTZU7
NGiWhJarGZj0FPB6zcgn9if3MFH0snbN1Xq7ZMaFsFgblc5eH/C/prmUqIHW/Amqk7lsAk5ScsY4
3HT3k8qMhEee+Elf+KRkQUUM7PqbNPogm7vaZLNUG1VSCe2ztTPfrOhw+rZFR80IE62zafLdOy4l
psQKeQq6cwk3fHHWBfV8X1qClgUwa2HB2towx/q2Xks0v/dkKwD0bR1w5YMHlesK/JpgQVPrbeN6
0VAqruXbBAyTHuCvZHZqK27SsUkrrheiFiBFJthEEYyJ4zLKFrpN5PcxZ4cK+FoyV4oIlQg3ocVh
+n/zq0vMMEMVGs+OM2yT1ugSsFHh8WrtPeABYlbOdTkOvKmyyUdsiIb3dtrF/1v5js33EAtGMnQ7
FoHZ/+kPIhLb5IIVPXNxMSAbjGnrCrI2Lcv+JvEbKfEeescCJqIOEIN2zZmu5O7sFz9+3UMjcCbY
TmhZANW1zgVTpdjJhK7lPm9AkgtqWV0Nl0q7yRewjmvMThGL7+L1dMDYh3Md42zQCkS1Og+P6qop
PZiyaCNJ1TfL9NXKMoFjAfzmXKKqBynZKxFFqpmFsMGTJZ/P6oWgioSo4bS4KVEHtpjUyiaj5c9J
e9TmqG3DUORHDsxXqLVe/kyM1yzZ9iGrTBrL2gzgy/Zwaet8g01WBdNCaLJEpq9NfI+r7EIhJOml
Ef8Y+yHGZfiBhx2mXKDU80hTe8Y5ztlgE3RKSOKjZukp2V5PoDzu+wo8iVF0gPQO+9jqR0lJIUtX
w7F/ZENWA/EYx5ldCXBYeVFX4kZLC8Yj40Z71vKxh4LF37HYH9VJfvlqPZ508vS8zCfbvvTmViim
tRvX33EKLb2WSvGsCmmvOGgPxmc8DF+ZV8XQV9dbg32hpuET89Txu6ru2TFLbIKzCfsSNMLHVrKi
whg3qXPuqPn8K8AukRyFiONBH40pNZZrLZjjfIintcy1zaoWi3T2cFZLNH74bCZe3Q1PtefwSYiE
bhDVbjKvUWlis9yVPmqXULZXxU25SjHq4g2gKAVrOQYhfZs6f34MPNe1qnUeyICLqTu/Y5dFckEt
JvhGhPB1ssHAnQoI5NOTnCKjMIJzeNwaOyS/GBr3/xYctYGCKSM5Q+/9guyjsSNlUfwYbD0ETFQE
O4Ne5jhZ3EVBwwaYis5cZQDWdRubCw0M9BlWasPoRhtdFIqWr/rcWGJSMJgz8fBKc2FTze6qEEj1
3l9TUfs6JJ/FeCesh6RbJ39Udt32Ce/I5BsM5cyZrDSBSTq6wn6LRh0wZ0hNcEuDYdw0V/Q+Zl76
xKwVDlNAloe/OhmfTgT2CTRpZdVI5NR9HnStfIBYRYEUVbnhzFlQYoNabtzLuWEI0U6hKATqCNXZ
Y2odncVHboTRe57j/zCbqmfAgdht6SL98LTc+HgvmkITOxH3qkHVTgxaIwRqK/rvHvXp0O/fs/bU
v/ByHq1Bs7AfWwYLN/xiqIfemMn80nikRWYkymWcsRT6fuh47aBPTlIdrem3wgVakRCxxx6XaX4a
gnNLYaO1CaZ48lxS2Oa94SIy1aWA/fW7DjW5XKiLikLm9hBMt3QpyH2v/1nZ7dqzVnoD/5ewON2C
ymVDZCBzmMbUfnSHOVAcdcQ54+bDB936COPldJk+VZD4mRl7PBdoTGAfNPgwuQ9L3ipTF0eZau6r
Lc6qtBoQmYaEbbSKqO+E+oSudDnSi6keKCrkVCoabFaz/JdHixlcT8MWPbolrUp+7z4YiJrCSwnJ
k8cxvUvQU3DXIGVVwOlLeMTdK4pSsjmBXXVO3mstZFrr6rwAx6lPcnjJdjiOQEb2enRls1/dW32q
iva6EGWrwEJB6MlYL8yoLydr6XW/TqIveZA7tEQdJSvCGVoPupFmhtqcc7xOc7/5i4OIdJF7QtXm
ChxZsr6wGocC0+E0TrgelyDquT9pOSVBc5G17nKjHA/VMBlZtpugDTamNEdxqbt+bykF3krIGxlr
ou1AlJH9a7mOkCZtMDO4rykV4aWN+3ROO69IY8BT5qUA0lXbodU2zEgqZnu7ETpDThw+vlSamBtO
YLrgcaraU0u5qALu3ebqc76MQTHLgbaFPrUhICzeY+YitrJ93gUM37dY8vHJfRyFE1qxZACl3tB6
SWI7Nuqicfp0gQWAwlKtnPoHdoFIeGWpv1FiWzmWfb0EDuDD+cQJNDdBWmUQVVYJ1TM/HP7NvPfH
3FJj8XBmWRHZzJebxjCfr3PT30hePSWsUDkgzaUp2eFY/EATHejJtelpsQQy78Whtv2kxVNnmS/7
P98oQRAG94zMZ/iccocxqqpVfnSYes6fwuG8QK9F1DB90mWQjtpBxcGofEzNYnSXtM2SI/ghCNrv
iYQeKx48NkUf86OXeDnMyw4dRVjGbXNqo6aEiJld62PYzRzHuSOVb8Q7nK/lkk+4pUKqAkbU2LZj
9B7B1Ki4jRSKdMMcXQRKcGJ2IJ0ANXcxYnUJEyPxR6sZ9ry18CK1383AgYRP/pWddqewB1x64aMA
fU7kWoO5K9vdKMpVNqy1WXUWpq3cf5Udk8M/mEu5fgz5K+sLXWkrhfghG0gNahUHhebwM4TYoXj8
6TrlXQqVxipv7VcGeZVxYApx979wHApkuZuVS3qQapSjajXFC220N8SRCF+fZbZOf1+1afmGnLeF
jShEZGWepa3UbE+ZFO75rqP0/NpvOfsb0ge/7Qx99QL4kFe852kWYKemRXk7u7vab8600BXLzg+t
/u7t+mNqrU4F6CSTFNCgGIkDARB3+1RF8vG0Ck4CJHHYn6/n+bKkblQYps8csnhwCc9kr90xPBuI
QM0TCX63xDkY97bM2wOf1lD8cvdhGkG40AgpTu4gxkzl3ONGdNcOfFtL21gblqORLTmLivmnk+o+
3idoeeMtGChXU4y2tl5CJfi4vfbfQ0DqtoIk3/88P14FtWCCnK4LGYugXJZV9GMqGMCpMmp4k/TD
/ogEYcfANCRcUPUUvQB56MmPF7/THCfGW9NfS6L/lwtPe/cgFr0iNGFBPaa5N9nPSQJt60PWPCac
PW4WnABb5EVpuZh9vOnNNGmhx4u+21TWfUXUbL4LWNRVAe7aNyk4z3uoRA8DtygJJfpmSqd8zvmn
zYzwhkDlKmV+wg2D3VNalgs+6X9lS000I0+KsRGAu/ExtW//xkByzEjqwksgKtp495xnaPmr3Mj7
kFF3KscxQjIMAqlhbSz9P9Ge4C48SfQxUnSc6cGN1urVeA7JMYHDN3knYFvxyAnPEkfWUZlCK4CO
IJvlDNcxQiiq2i0WHoXQVj6a8DT0leXQjrccvvnWRCYdYja6WTgbJHb6w8+lHJbaiWeBfveGPa0Z
nXCjTPWKEAvTlnoRYWj5LWM01OeJRjJ38o+o15W+HjfxbuQeBJ1XoFFewcrdVpF/DQzqy+r2WSG2
tIO5WJb9fNhOdEmpFvs+7RTMwAXf1s2OIjLCIYsjjnBM7DxdwgUYFj4txEjLICRUoSO7S0Lsupx8
E/KgGE91lmK4Z2Nm+hPesBcuTojq5Y7jZIDDscrUERROP0B3M2RwYjWAknmHPW7E+QYI9vzOUz92
/dFy+54y131msN7qtCcSxnap1cn68tidmVkm8DvK2B1AZ0KTiwQkolPZ8wE18yy60xZOacjiUZY7
bjMOBmH583GDKEoMLT+kj9XJ6LrxTOEJlYm2aL4zyoeQoqFqFGLkSDiaenrjt+29zZckFw+j0UYt
WXDtpfSlfa+Mu2SsdwrMj+tIktaFF/q0fShUAp2puGH3iqmzQpccGSTOCZi20JKRtJjJsZ+HwfA1
0zc2hT6SoqAVG6N55w3wvMTVatlGO+4DYHCml1pG3a5sAXim+LHz6PKw/QYGFylURHRm7/I+LOTe
663KWqzzCZ1NoI7Xpk1g8yiY5JwoHfv7y2SAX2Zh+RHbLieKgKYT5zKb6ionTzNyb4BLQzePQkTy
DPBCUQ8jTrWjY0OHcpg/LJiPPo2nd6Xv7Zr+N5PyqOG7XtL+A7VRSOkSigThBVfjQ9mcpUGEowyh
fS2jxgc7oF7QRJsmCcn5Ebqg9AibV5URbqsuMTuhymmtF+nPTL9dy651/ZBcl0/CTcYnU5thdMkL
nx+sUBScvNwZ9+ixRI3+wxhcQ/r4JQ6xcMeR39ZYupjI1+btFqYxr+M8NyWboA2+7uE7DD+HdORJ
32ExPJVzMezxns8T4TAKpy21CyHRbevi1SeZyUxVL2Gd3r+TcvBWDzx7fX3B9+oDSQN6u7Q5aF0A
Wg9hLzURYQlt5Szo5so9CMSg8bjr5zCL939r/nXDdgJJcddewOwPMWxI/xhKYB+h0cxOv5/E2vn9
7c6eJzcCGgKxc/3axUMF8ANy832xE7Lylo8qnX2+cMPOS9atwu0zBsSlbdx0G2QoV7KWoNYAIsMp
FQuPFyGjXFSvSvjNcg2rxGWmSsEMFFFTyHlVqZL1++cqaGkoKYXQX0ymRpDYxK5+A6+a78OFIu2q
v6zDFZLSVgvQ589cdB2o8rcOrwRTsgFfrnF8RfKcyLiWm8QPRCOK/N80JXSvh+VriFTsdkcSvEhW
5lQScQ4mkJiVIYeqfCNZWNnOqy/eM6ezJFzvdisf4Qc7XKtNKW/rhSHxDPviKcUQM8dRqf1Kdhc/
BjO3wdSfQAIRS/IRryUZC5HTlj1CEb6JiKxLn+v1Oouy87/AUOO7ZtmNJyr3B327ChwC2/8TWAt4
lw6XNEd3PFgguqZ1i5YWYdws7euB6RIeSvncJAEYA3RjzH+VCvDH//ZvFDvwHNtr8h9CKGNkmYO0
AbzG06lLJIQdj+/k7lnRatUbE2eQ/zYpOINq5LuDgs52q8ss2sMnFsq9W5xDldwHYfxjKfSI94ma
/ICVYX+B2yHH0D60kQWsHomEo7RKaNC+gM66LtBU4aVWsXISWSujCLACx/XszIVobLW3kKd9XbUT
jj4tedUZ3r9c9s2AmDlndMtJUydGfCFIS9p7kRsJSYM9gfVfeZL5Ma7taFovdbLTFyxskDT0lyuU
gBvQGc8IpQXVYa+EH1Qcsbn19//Z64DqV5jZk3d19mAMKtAD570B5iVeUaQLj2b9DegN9QEd7v3I
mfNbIAi4CyuGQjvznBnlykhH8qVlQATWd8KQawuQcfq5h1/2JeN7Fo9WQbyS/XC9imIAPrFU3ROK
YFqmSGdZmpjHkGcc/Icc+7nEj492c0HtZ4YKNSYfdrwZDdqZcCBKkE0kyCdRF0MCq+fCRPOmlkZW
CkszbmFk54voo2t6a4wM5JAOh/v2cXqmA/gbNe3WBOBCOKAdMw2apKUWy13gBrxXlbMpoPgh1vIM
MyRX9+Td0dNrVEUkOWiuWHyMeiWqHTt5O60WVJY7AGG5fJTimhVFQM8uizVW8IV7JzxKESfbCS5R
mvaOv4kDnhiQP8VbPM3Xv7cxcoVXRaaYpbsCS4TAaMOOnCcQ0V0duJKS0I5+xF2/qZCqSJmjYrXC
amsagWQO75fctE1FlyQVgVpmqXJH/NiSgDUFhULV/JseO9yNfDo9xS0tP7YxYMoucfzW5ipYqcgU
BHHrj+67k/pjTXCfAocvOD0BI6E+qQHHbn02i05fQc3lvsHF3Gw5y/lGdn+RulTtf/ikbAlnCcgy
P/gAvCdROKwThVP2PV4WXWsVLjWHau8+nMkRPo+d5egfGLFFJEQcrLEkEJZ8GQkM3i//AXmRXdLd
10s1JpxYb6y602TgMz/Gnn2/VEalPUShyKbd9e+/h5kdxYfcO1gSLkz9d0QxkGJsXHqmq3R1YZOo
/w/903Yrdam80ABCg85/j6OrSVN7dmysUf1rwUMnikBeyoQAOO8PmE64o8kk827opj45WVhhYqZI
Tpl4lx6xAMsRY/rDzHeg0jZYslG4QtT6wwIt6kJrI0bJU/eA+A95JuGYYqX9GfKTVIM2LfVY+Idx
uoJXP5RZU1jJGBSiFuD00UIpUUVWAxWNnZPx0zwpgnwDuOjLcwyELVsUAlQm244+LHZEYak7g/yS
BVwqubCtxMfS9MINu18J8hSXWEqCuJL4BqJgFtdF+GoYmUmx50pbNSPta2Uf6ref+oTmdud5bTIN
uvuiR/vv4m2CHw9NnD/aobujb1Rp/wGGEr7NIT+gEH/awaKWe4Rtbp0UNsBjT420zEZn1y4ByB5U
8GzcRYAMFAk+qrnOy6ga81OAdQpszDKAwO1iSGhjVaOss4kg54j7tTTP8YygbSAlXEHJD73NSCV0
w5Dldfwi+d6ebQW6mGyDA2bZKs7W8Tb06wLps4drDtKsQjeUKNpzm9KtCCGqVcG62XNiqfePTrVA
lpbeW+6tD6dVqAx8WR2w39sdqWoX7Z0Ql9csOmLZJXE67r20vSerqAHo/mCgG2+DTSw+HFoV457e
HKSFPQ6YOnBI6gB3x5U8RdmkkF8eJeR0HvpGz7dmJ+u2/3gJ61tomjZoVATKEvmlVsqJpyq+SEaR
GDzxMQ1F42i84CXw+HxQebqz80C/fD5MX+xEUD+vCLT/he1KO/2IZ2mK8hSzH/iiu6PIPAi1NK9v
XEMM16TlrQV2nmczyiLMLT7uRoV2qU0gcS4v+nqnQ8goartbFNX/BG1T2qShVs4YCB+vt5PyLUXR
pm9P7kh8fVMAGb8NCTgMjjhW8roee3REVUEWBFy+N1mszFKF5ZiI7Llm+uWki494BdzEJXaJEql4
MCWlDbejKB5Z1ycvaLmb9s7KzSs3/M1E9iTVxZwFsiRxUwr0RW2JY3ym0vz50MvJzpWpe1+Q1jaG
uzuSEHxapKSqa2baIWgcqfwYZQOTdQseMnyWVW1NI/C1hyz7yjWKKA8bWxgGkpzp9g2AhI1jUISd
kYiLHrb81ehttZmixhKiGhq4A+7pOu/XzcSXt/DO8vq4fis471DfCaUV1YjZYp5meX/BdtlNiuy5
pGwtJeJ8HMpUiQbW2du+HLnTO8I2HfJ13lJWhLMneGq2PbaLK6gitPentR/26mx88BLugO+uH5F1
FLyZEkVgTTcZkFmQZRgjK/F4fKE1qabg7TPtiZ2zYnAjxHtuj0XaoET+xQmHsmg1A4oNmPQydFzi
aF+gFba63lws7dg6xKVUA2+Xl5wUj9DwLuMLflc2xLx6fG1XmV4S8hQQ4h5DU/StUeJ4EDc+F1mQ
Cyj+r8ML8n+ZAQveR3cQWgVX2vkMbBllsXXaTHwdSzTJqWk7L/Ud2nluRrZf/DOU0Jq7Q7nAczRI
ydPYAK33Im3S7qr8ZcFaykCtICU1XuI7oeHHGSSBt+00jyr4yHPOUMe3UdkknEltJi/5SCGqOy+F
TNQFdt+rP9D2lub9KZvxJ5IgZ1MUfoSnZH48/sgW+dW7d2qhH1cCqL+WlCMX3XSGynRiPsWjAI6G
fptDH3TNP8CJartwcObUrm92HBhbxJ01CyDXD/LKPJQs6YBixry42msPWJgeg1LC4lh35NViPNU3
Rx/UzRoMBsjWHuTLP8pkSUxdAamCFkErVt7f8/jUL6KcuyqAB0rHxyiPg9X1AkTRQ/BQmvgTpfz5
7wNOt7L6SndZSnelVBoQGeuHE8QzG+EL6zm9965aMLFmU29ge/pMZVi2b3rbJoP3dz8d0mh4spcu
5Ctja6VD0ZUaXG0I3/2gmySIalOYuVh2j3oBzD78mWkcbqKDMhIiCcV62uI6vOv9cgt4ZAX8+QRC
qSAVPxOeNItJyAizY4GQjB9bUxSPiqR4QkD0XXTiW08htKhZxig6Heol/nAHpocID0R2JvAYs2Vg
VeouRz+whtYEtmzHJ2oZ8qB1YlH/HOyD+2Z26dmQ3bg+zc2crHqxzwPed1nZ352+JTOEdCfv4X1n
ZF1oH5Oatv9d4QySxXUFSSZqJSBDEVLRVENj+8+03rp494qTKlpAnvvBprXQYaYrxXt7HAZe5nTi
b2I3/7jznDVTJ+GEnSFmasgf5U+a3ChqvLEQQj50Y9bBmZtTieZUBilokDuIv61DqTHiJC6cuJEg
ahcMIKonKHklF7Rb0PAosOcZQ8sQ6l4h5U15W9SYjDyUfFaq4ZTH/f9hWdekrMKQUP3bCqqQNM+w
Uo4wUVfGOhRTRu8QXNElJbk+eFIvuF1aLiIT2OLfP5rbFSiHH8w/ihCcLx6ctUnf0EqmB0O/KYio
sWDyLBxsX/abITffNop1iIQjWUBE6/zfG6t373v+m9x0r/bS+TSmnNFgU6xQfXoBHsg/S0cKi29L
tljsnyK4i2N08w4E5lZBeomWZzZNFhxPoMI7fktdPzkqy5oweCJhHUiYVaOm+lHNtzKKV01UxBGw
0PmhSEQorW9utbvpJZxDbg3TmhtlZK0Egy5Z3UhuK61wuE4kmcMYUHjRDG0J/A2WM3KvwI85RVIp
6iQr9xTQjcCUt3eS4jlR6v5oCnCPv5CJKsZpGO3c8I3YCGSOC+xB2df8wFM0fJluy9KGaPedrv1+
jfQRlLj8KSPA2eB5XqB8BBcEoH1FpKqVAvL3S4LPALA7QEcOAiRHbWPs/fCt/9/g+87iCm1t6CQQ
A+LmP9fD6x2JdbGOYKdZncMqFUeDA0P5Wt/7KJ+C74I1HmKJAApBepJaS/4eZrYTlYfuV/BjJG0Z
dYalJYLEDjOWnA4Kn4SEx07s/rZPiJ7bBOB0gau80TcEyPvkt3S5NRGFA4NrymwAvvq0tqeqJ3Wg
+sGvOzeWfiPLtVEbxhTYF1Sh1iCL4t+w5ZFDixn9NhN3OOpczDXe4+SfDFIgfDIAs2r0+2qi2yb6
XuGcyAcTYQGxNoIUcCMAz+XLEVjWyujfMsg8l8pxEKjCXkaC0/kw+VP3GGzCWRqhBTQ1LTp5F38i
YrXj//QJoCvPrn47ufL8gBWWUqMK70WiggAa3Wb2uaDMmDhRsOXVBTFFsS1t3nKxCC+mrKslP+yr
OEqiZH7uBTsWGl6X+qE2dNR/B6lvIbcG47WikmqYeEPZWxHSG/gGi9/pAShzbUvWWRnn0CnMTyub
dtlL1bsLlAMY54tk+rnYCbY9DH7BIIbvbXeKADV9MVM/VNN0dDP1Wu5yFxJweoHzUL/fzH4rMcAz
NaUW/GtM6mym05hT/tgHW60Nu161MelasB0zbS69xRuOM6QJ39pxRGZ1aeDLxsB/FSfwzBQQydZp
UqEededGixQIXFDaZk3wbuISzrXFD2AgiLQ+jL6jHAmV9FwMhMKnLHHzLhliP2dngLgQzm+0g0qS
RGiIk8IIzn9lq+ZYVigLxlnQIZzZlbYu3q9KIPmvBdkduENwmOi3/CprBBHNRx6T/RaaD1NPyQb/
q8sKgNy7KDREbWPdNwa50XwtG1NZnF/rxxSOuC6lsQywDLKSur4LUJbIolDpKV43au9xobjvkRxL
0W7p/MvXFSvzdoPu7FpS0Krr9XHoo7ve8fazcRvlQduso9R9cwsBc1r0TGK+TKAZnOoPlfAvoO0V
GNzh6iRjiq2JNUIkAmiYNxyLWMmVg8e8So2WZLd7axVB4/kNOWgMRVvXXukXHK5RAXYhv1KZJ9sC
zBCJlb6DMMoU/B2aiUzBfkaWybh4JSq6EiJ05gmZfU+5sfWO29wzVVwLcleIDjHicwyZl5ciLWEE
NhK9oWZ2UlKvAHed0eiI5uMj1BQARnQaZ6R2a0hUZ48hsEyPlsOtkak3tuPQxoqPSY11Gb2Dvjyu
kR0u4UHkg8Z1QezKpXQmHNSu0Zc5WU4g27wOdiv1HKRolFFHRyvnBOtLayGd5bb5po/7VTRkyqYq
2q7WtYGjGj9QA8PUSPv17UVTVEc/zLtj0puymd/IwVB/eMQd6gDZk9m0cR7+yXzRhUk6Eq/OE+R0
kmtgAurl4mVBw65kfrGzbSPQa/mVsJqgh2j5vp6s1VQIxNQtJKGYMdBJywjypjL/nG44ZzoX5F1c
/tozatC09cBXnoaF4g4a9NHGCfpT0D4xksm96a++u+v6P/fTW3iMeJjfNalzqTnwNJcZhkhz9wj0
bLmYYbukpQ8QumtRn7lStWxooDej4+lEVks8vvhdri2jHb9WlfIjR7dWGN/+pSyrRDiTP632kxed
DR00JMfwvsH4TqPBRz4hjfWcrUVrnilmQhxxXRjCyl1lHINvdKOJr08cnXF2YSBYAxHKfYsbPSTd
aknU2rvuiKMhBY7qVQMfVhZZnZWBdSpGYHMFIfJSCaKGY/3fkdJyUjl164c7ArTMx3vgq32RAysw
sVmK0ACNU44NxZzolM66ZOSBO0XXq41lJEK0KUWUS0he7muPsYU6gTVkeZn6Q23BMswNr0wrUhnD
kiWDBWZ3vxy+A5qbOgwmgP6Hy8Sj1ICIeM2rsT9qRwJl6dbmm470ADEvh5IHRfesJE16SdElOV1m
nrCYZc5csoUUgkMujuFOE1Hscgv+uYzduIKUwIGbtKmaDGTw4VzEN1pF5cENIYpZq/x7ZSfaVbKu
C8sY9zp/jZkLWp73pVawQaKNEMY4LIurOHneP0ZFnt1abvEfdHC9+RFJLfQJG56AHZNnBKnVtZ+e
/IumUk03hYNO8zrHX+1NT5G/+ClG1NtNQ1JATVkm3u3u/EDGwPH67O0NqWvBtvWPBEwsMLgY5XLB
xBGEivKhgfzcrXjUhKgAzVg1uAWAkipc/wCRjrPRBXtROJerJvy8sapqgkwbXN2dceE0rTIND7Ey
1iMjpEur0D3yZgLR87/IfoE90UpLwqJe6em2xKKBTW4YNwPhHG1NMEVXZbpp3i1p1tW1SUaAtfqU
WVmWmalBNcdFdZAYUaU4zbbjIBF6RLvZ7kD5PiEtTY9CpbPSfllsrvsBpdiVy9FrJSfeDxr5GK8g
Si301M0Cym0g7fFDq+gy/MZCgnDwQEc42+lfmT7qQru2Nd8B9OEHK0uCEYq43V5wxzD1OQ/gMP15
7v9pos1beR2cR8Lf4pdFNn8rZB7aTpBwclUykxQ5XmLrhmyQKDOjyBi5Ulr4jgT3f8CBg4+4SW92
yuA6pz15DJT23vZ5LFEAbvM8HC0Isv+4Lj0n0fQrRPNBVOE7kzqLVim/zkJPZiibR/1SBtT/RHKG
nUuW4ZsEcEh5h2Gd3NplkGNd+hjU/EFPChgu+5DaagZGtPzSwzRyxwVXtev2V2fmPK9P2KOU2E1I
zrij+JlE2JWIKWPRBWY5np0f2GBE1JGNVt2TfD/LhUJqeqUg1g5K6UMI0zrL6jCYgqTJXLlIULu2
txnA/6a0JOuvdPv4mlpThuxusn1Q2Mi4Mj6d6MF2UL89Y26brhaUyZsu1UiDqH5rmYgH2aNjq7g3
DvKp93XYrHj6zir6PHKEX++xkqpACrHdKIxkZ51oFcyw+hHnySTlXe3aZhFlAuFHQBmIEwKQHAsE
mwdAyQOf29EUuplM0hnHDGmBC0ijJQpcoRJbsSyaHPhWClu8QDgA7s8cxb+bTwrQAk+t/BT+YaWI
HFgWzCbMooh4Eecoo4XWKdQwoOFHteBXPObo+FB6C2mV0q04TzChBahE8dghvlemhEmvuAnGH/um
9BVG8lGJQfhdlWwIr3MRkJUZuJ/CFBf0XmBTcdR+a2u3Hb2CbzQZPLsOnb9f2Eou8vuod4HYUMV2
LMKZKvGQ+VASOfULvO6nt9x4khmShBRZOSGJcsqgkkjnY8fnhAWe0akCchKS2oByTC00sxLUei1o
ES6wd8aAax9+0kL40EDThRJNgd0AimcnoEaNOeeT3oNWku5fDGs77mxEnVeM4NdL2nACcCipK81o
GwRrIWq+s+0WfraZJsNA9RwuWzkBOXp6Dc4sJbk3U76UIEeBLmFZUBDy5d6niF418lru5bLWQr5U
dgXurBGU5wzOITM6GRMJpWx6JiDZ7vME48pmnyh8QxRH6S45YPYFfPRTMd/2KWuyXbkUvB1vHpnk
G1Cqx4mc6aF0dtI98xI5/89hOi+wfDEYmf5KUoneMz8oE8os05L7Z9TuR1FCj8wU1PwuorpEaf4x
OjphDGictyJsu3pyc3Jbki2AiirNExgiNLoWv+7lxCMrxnTm864CZ0IDLRhme8VakmSW26vVckRF
+UwUnokwroxYvE7M6LBgV/xO/fvb9pHP+1Bw/0w6TE2RtkIsqaYudwwESmnPLIziGD7kS0hyIIUW
T93N0WUQWbztgMVY3/z6MzEMCTPD85HGpaLfxPFMfnkgk8x/W8elqIf5i6IXEhfwnx9cn+EaIWyj
SilRUAoDQBvfGQeS6/mShgmaG+t655ux3Gl+HjVZ+Nbfc1k0gUE0KIDJsLJQtVp9m9mpBQUekrnS
uGthJqMgMaTzeqC/kBchChwLb+C31ri/a0Zs+jXhkAeAO+6SEKIstaSPMdOO65JBlv9qNMha8n/h
iBiHwx/S3U6NuEUIzSRlv4r1AFtnFKjKnULzp44ZwLJNtkxrWCkXqGw+uPmByfd7FxCKypNXdNfo
ecMyhXIvi7hi2K9wo3dLrq1l0YdcC+AymFvgGYgP7u6/paSG9Jt9PA4vB2/I38OSM3kQ07wbpKJE
uQ3momJEGSHTjSHSbRtALkoXUcWKMu18yd5qmRGMJ3/T6WAgz+UJVXpVrp09Hu64U9BKt+gfKJ9O
1g0AyAmg/eqGalo+G+aR62yQ29j8EnYDSMCeSRsTw82WYO9aEY+Ep+dbx2XcrA/dnSJxYXfH9VWf
TlCQWMm6uS0Uv4JkCkQu61lKqaX+2iNhTKczuCqgoiymsYsS0SOJJnKt3dHlKzERlmKCdqfeJciq
Ceo1ieHQkT/R0kV4YmxKxw2CjvcLhQ8BFoY4GaASQj7DcFE7Q9Ch6j9+X/4EOE5blDlHnILxh+o7
VFgI8dxGFVKS7lgrnszJDR0qL2sui8ioAc1GT6Kd+X4ykCrRc95J3R7g4MfLBE35lLFuapyADFSN
zMSPsLjnZTC+yvLavjdCWCQZH6IqbrrI1kmcxFvq9L6ThMrcW1jQPteFFx3Gijm7+ChbtH2MRYex
T+b5gBu50QYzZoF2c1rzT1XFyJS2b9hyPN6WBQarApX/+Kr0uAlOuh+3Z7lKCZrQCj7MfyJ2WNIv
qf2PY9/4TyfoeiBQKC6iWKeiCWp85V9tjRTBOfxSwLnYU5f0F0m3k4zepLt/ZbwMK5fWFuV8QUj+
Uy9TN4x8S82zpm31kpLL4t1KfDHTSo59pO0SW34wBlK1mOiUjSfSWuGYALrVSebdXADJkKHlbxYQ
AjxeDuQ5Oil5eA/PmB7AIb+5x4vvyZ5Qkx7WXYqrFgduNdGLqNYN8/AEYF0di1imqZdB+Irhl2qp
upbEDbx+oDCrjZ5AFS2FyXbfZR+2XWJrBiCzBLVVb026WojbGjbK5woDLYD7PLPA4maWsXCBfbin
J9vGAnwQHEdcLAKku9XtUO51SWI0BAUMDaWdzSsmQxi0Y2bxF3veX/7SdpCeCJ8q0TQ/tOk2Vhjw
OO0PlvYSj2v19M9NlbofeWXnECiaHmcC+8TGp4cmfNoideINrTi3D9QuNF9VVJsQDsH8RZwAdibE
k52a5pjnofUzEtR0KEFzrcS+Z7qzqYWFP2WR5f3YCVG9uDtp7JAjOD/PbiD5uXN0w68Cds3+njYx
no65NSzFaQwNMxCRipbx4QKHie4ExiC8rnTBqNzVLTvN3NNXEL3crd7pGCBbBdMkd247U4PWbnhB
8D0qPHRfC3hXZyibU/W8MmqMpe+kmylwerv8/IfH3z8q4lX/QTwN2gWQMohvnXAxhnEMsBPp5bMQ
GwvyEIu4uw+foQnFZ4GI5x+Je4T9HsuhTR+AChKkRHiVz58dOhkP0aCQ1Y1zx3Jnuk8fJRBd4dyM
VWMvS6iSrjmV6xkYDzJMtrBqr5jzeVwCl1+OFqHQSNgIvWvnwc5ybaImQZ3sPj4wX8Tue1Z0P/QP
Veq5fJkHo1sW5dffPhXCt26RORpH5R/r0z9GOlyh7s5iL+iBRL4DwOFJCKr0J1F9ypdmpvioxWcZ
VQGPuU4VviW0MSqbAgIJJU9FjQwB89FYezsu9fbsh3TwRX3J0H6BZIGgDm0wOcmhbTW7ZBJLO0dt
/dDv9EEBgJQVztxgrzXgv6gaYqWINHoEMeqmPPgfnwxhi+8wFEfpgYB6FrmfhSfYGD6p7FEzr8OL
GezJlVLh6nc/yY7m56NEY2RlUSxgUPd/J088Bso8oyipBhgZ+vaY31+j/7/ItHBiLp+y9yCbfg7W
oyy6l6oKVwAFCJUoFUAvxRlzHDdTT04ChdX6IZ0RspS3XNzol0RsXhtYPI4KtRnafsHwvkTbh7ok
mCiAm3dZXS/S9hPtKRFgw5AsHsd952Yanjeoracumk1wmFl7210CqB8DHAYS7/uO23eojfqmPuNQ
ky9GB4rkCmIIfZTNK3ok/+9WlNMyt3OVAZrzDa6AmEB8JO42c4S4GV0UW8a9ASsJaPFZbXycIoKN
SK7DW6qNQO75svC02fv8f5ir+m4enRFX8oiWcO2pEOOLLNzrcEjMn0j8eME2E4xIxwxEky2WFdIi
szFwE7sOqwFZMD3eCf9nENszMinskbw8ZeRQRIjw8kN54S9gWt9F5XvddcAH8OJ6cz6UaQdHMJN9
UBRqCW2A9UQLl9goKDlXa9QHB3HgrCFf5IXVZCz2t7KbYMsJ/LmiRsPMksCulhMg9rWrleVlam3+
i1cwLtrczrPGFGBNB9qTveElWnPwoEgiroNkG0s7DBpJ+uFpHK5HCKuQrAqT19BAjzjLBz2jTqMx
FvtsQFmZedUiEKwVoaJk0tbEyaX2I4LcR1WJfwHg7O/Eq7t897uLLtjGPz70Gb+GCQ13+SGb4dtg
IHlJTCWSNMAvumPUZ+8uwNtfDIbCLSRkw9ZSh0P1BxPsUhKedspP9Vh+/BkMsKEQFiRhnoejQf4I
9C+qBayV6ephbtP8rI7gwSLYrjeybLHi1dHYleTk8fWViiBn2TfEq7egFxkDLHJ3sH69r8MOqvok
zF6our5XTtdIdVI2qFP4dBDPQFSMsELLlvpL57GycApOH1h41lgmnNiWs80VDD+QK2lcimKQlmKr
dRUH6NA3KGVvXhMBzoozAExdGkohVoc6q4PP6/p2xfXPriB/cGg2DVsFZmmTYGOOHIe8vPJQsjhK
EjMAD1+4EQnrhN23yqFCEisI9o469/iZyoUl01THe32vjwKlJX2DG5FCzpc5xRhri6V6r7i+qe3G
ZMCkmev1SLoj1TyDRtKExYShAW7WxuBZ0Gbt/r8a5lPxrcHh/nelqApsXZQGISeb4AZMB4/rIqTW
f6PXCykrEoITo+kyMxgzXIquk9EAewmaqJ+DE8ugzgDStSNwK5CaXfn4VTooGrinMsbJ2xFklo/X
q9EyD6vhDfQlXEfe4kxyx2LMsVpNFwWSbJaywl8iNUTTo+SjVIDy54jdPtlPtxumb8Gmt2jmLiEh
27MC2Ykqvnkf2iFUUYrDo90ijRH26zC+sbeSzRa7FOlFB4wMM2JEnyLFzxN/lUCKwu/k/jUy0RjT
RAK864h6ucr2myc/IqFDdE7MNKozwpBsRKmdJ8MqZFuzWkaY7KzoeTTqYzVQxoA1Ejx+JtCpaSrx
I/wBLmkQIUqHNDTQSAshfw8BGaRuIAvOa0LWsQZeqoUYm3DT5KvS8aSQ2E7n223h4pVVFM/MQfXX
KY+/urgW00ONZQ+w6puC9ZxqqqLWo5xhxSOM+RivMXDxWgFElVoU4WDa0RUSWM9peV7J+17vUffS
m8M1LxMd0Nfsqrtw44xnoaIatNybwCbBK3h8n3ToOjVLK794miRDVNG8AB+DM5jsJOs7Nsk9FASL
dE97HNXuQBz2t2nup55KWRMqt+oiAGUfRoIxOY8S3nMk7IvFwOfCujXEp8TITX1IrU4gugRttNkB
ZIG/v92UmGb9FGGdaEAPUEOjdhJCfy2oTBEnaWX4iSpZdfae6S/YtR4mREOeYtId6PxAPlpcFO+p
TEnuyOsOfTHdZQ0lGITHUEHCeoAwygYhf5i4pJqLvbmu6+fGIEIJ2xppVrFsvhPGG/qMsATc66Zm
bkyfiRdKbSQCCZZFrQu/Tn1JOTsxIGo1eqvpcb9Be4uOleRfk4ON9pPVn29aoOC5KmY9t9qgfDUf
e13Jhcs3+ADSunH03UEAwmGgMgkiMjdUR5ES6vr50fc8HHpfN1mpJTSkzaIlB9LwpWkAg7KVJ3Ku
YxYmD2lQrXVcE22LKOMWcmFBOf3iVmvY5J/JFT7JNkxpB5eHAVhCFPhXyNnLfYbXoirdCfq54k9F
P4NefswieqA/3/2s3fF8CYJFRnYvZFD7WD1FiZf35dI55hOaH4ErpfP4W0imOVh17hpVZXfDf3Xm
6bHpYp/sFTA3grD24hW2NO7MWxvHUmuakDMtTbV8B8aL5cs+/iyeiwdt+3CwI7zh+9ia+Mq7uyVa
HHsukPaPG35+L0KvsuOkfvqcOCBMh/TkpuCKnPU4y6h8b8wbB5dhAwwVJ7lGOCnE+LudrqKzwuWU
JKfAma7gfoWoENVDoICffC9qRRZwgCpLN+LW7dLIrcN6kb11R7ukvnTD2P5owMcKQ1H78vQqhnYf
UnI5FBUUrmv/94nxD55+8GVvih7fQnpG13hq8+kw9bYVBS77DgnDgKtutGqYG9pxrRrl8mU4v6sn
l7rSNT6Vyk6EkPUDToyQTZ5r7aP6oGhZHD9Xq9h9OihE1DZ5OlaX0oMQb+yD4IodKy5YcVR6IAPe
D6CmQfYGa+q/nZCpncazk0pzoPx8/St3rsZqgGqoVP6wb2ofgGUzkcX/H0YPcXuzFTooqASaVfer
RO2oe+rJqGEfic/TBH3fpkXxQIclFupDzPmlWyeMzv4voCnYTBTOHiVcx8rlJqDWxkwfS5UJwjBx
Ynef/paXe2pczmBMAaEbewZeLQvBRrYeDA9vZnYpa7jTEdu3yOXlL5QuZP84lcIiNhAiyiH5BS27
d5eXw4Gere1XiTM7Od9Hpp72QnG4JQ3GmFLYPHOfl9ID/Iz6E13FWr3eN30d6qkS7GY5n6DEzdCU
dIcYZHBSe380UxtWFhU6w7kHuk5i1CvUVzj0TqGAGavT3Mnta94RlxZa/2x3xyJNF+nqhcrUpnLK
Un4lwXoNM6M6yr4mIfWdFQKHtnrfawEqiQVmtxtyySpFDY7z9xAy9VN2+IK+Afybcdz19jfSsDih
5VgkViNdNz67bZOGX/n7CBh89ksq8fVewdNpAP6P7sKrdWoncQBqtPULy0FiaVvApcCTIKE71oAo
3sbYnsGiehckOCQpwylXFjjzP+LZ4b7mglyma0VtitLXFuFlNofqx3qpVsiWyX+yV83PNnXYSG26
u1HIKF551H7mm5uH/imvwZFcyfYimQ9GohhmXA2D7ALgrimGIgL2SRufw8H1Tn2bdwKN09EjoNwi
/CT4eV0TJm5e3yqtLFvqFNckxA9AFMiiQN2GZzlL0IB/zXgrLE6Vv1e/WB6UWqK2EjT1Dj/Hklln
l6vBNQKB2a1EfgSb9upCtX4cQgBmbiTSGDRwBIbFA4VTTbAFTy1afQTfteji/1ad0s4hXI4lTTiw
f9A9cwWiDS/mT9yjvnyzmA3Ah7SqZ9Of3LBkug2KRTg+RnKAKUnWKOn6llnmFGB2L+JIvT3zvpxw
qeyw0BYWXf98piNZ/SCP+/Kaa3q+yvaWjDL5Mautf5kyzRg/fKNk5cvMhA8wLWaFOOwZlcJx0UV0
2RSDtcPEkMZ1Zbyfff//3bqPqHr2zWD5QgnHIbR2h7pX2CyampNdH0AJesZSoGb4aHpvR61vv5bH
SRWam7kPA6WMglJkV6cGSCzVxJ7jcpbZlDfbBsoz+SqZEcJlMCq5nVncJy1Uk4kwSBZUwucN0f3V
mYbPqUqEVFFf8yxYPxSC9NGDWxd8twv0Qx8GhgjWEEEueKzSdp5VA/NzRyEZhsklOCzBXY+KukAV
9rO6COVkKFR+zRVD9rPFUmiY4qMrZXMuo/0Wj5sNuAwqy2bAIkv+VDOIvjj95kLWeEV5y1zFT8Yb
1YKGWv6jwWP42d3q7N/QcQHfCLle/4JuQbmWlop6sCU1H8Nq3uqC3v1ExyC14aFqLQT2GZ0mpPFu
5pT7uabfZtG8ikyVbmtvHIHioFnBIJ0fX0sguEIrJoOq1pcIuYgtJT/RzzWFMaLHLZI2cwqgMD5+
ZsYx1KHiyadCE3/MJcu5D6FhY5eTC1xJQU7At8p7QqkyxQLRCe4179WULppU4W+4HZf7h87SpL0M
jp2TE2yqTi384iZ6a0iaxG4I7QrJE09Bx0nEOwn/0wMc21esKZvihGWASNyyXSlNsehJKs3ErvvL
N9IKfFMRUxd17VMG1XdS7d/n72EvZ395OFJZxmlHebVGsao9WxU+IvRpuDdSPjM/jEOiKA9AE4gZ
+ogGX0PunlQo5yNJqR3/zjrbvanUYLsZs2Z4udg6XWb3AVopUtXqCpLh1jfMpzvkSAwlfDmcIbzV
a4j4Aug+Ch+gl6Vni/nyudn+xrNQT6YfO5ih7eLVbGnDTNCHrk+o8fTrdFnAyJ3BMhm6rq06BwHy
y2Zdu42oKi44oFXz0Zwce0ErPbZOCAJsoUGp/9HheHqeiCNCc2WvaLxxM9sVV2Exz+2ENY0t0USO
3VjXHKGGhh+8a67t6S4SsxmtVoKrHhubdG7RE+Gs/c8fCCNDrjr46dQqt0smfTy7tLBcKhtX/IeA
ltuorrpuhada4Xrk/+miMi1WTQ7szFW/wK+yuZ/NZtC+n5wprsDFh852O7nhzQS4h7umMQg7zYw+
lToKGpGZDwRANecLZJawscqrtpUqzrv07XRUn2hRSDJNuCVgz4rp0UdNHPbNm24a/KrPwmf0x1fV
aIstWUzMRIxezuxwlkS/7rLrWJ+NyWDTYOT8ypCx6w5vWXdllTYjIx5W+QmcCuXHzTpiI+9nqBl1
p7mCjhnvDr+IYogt6nqM3zmtnL5jVNsfe2QQG9IReCjqHkJKzxC1B8RxVnl4KBJduEx6fYDXUaxL
eLq8igZgnRDvw9Q98wEtg6l8mLYs+rpzazgCfko5KnbXdrBSs0R0Fv4YF4Qo0TkpILtvSpGiL4mj
MkL6RN7IwGqqffGgosZjbhxkxWNKknWu2jYnAxpb2+h1S5srbc3xBhwyMJL8ErkmtHSQVb1OGFEE
uKFi9pwbQb8qWFXco1COvUEJMNUh4aV4Qd66N3Of1SwKUXYT8f6OR3C7FjLRYQe/qIOlygQ3KNTM
ntVs9TAsbZ8KOFTvxHFbOmSjUD4his9DSUnqED0ZWfkCcoWkhuPx9wZZpXkSTJK+gbr2mfIBi8y/
no9LkMEDe6qJSnyNKQjGHIR3W1xpSDd/h6zVmUVDiopkUiM5kMRhQv609mM8cZ1+4pftXubH66/r
NhaixkbNkXMCFyZ7Bg6mXsB/3DKMg/wV38Xqp7/o9f26c/aOJ6G8cEWSiFfGiK5JGSl03wGUgtEz
akU62h2kTT9cC0DMGxLbnSs09BsEENZ5c9/GVASANZQL/ngbdLjg0dsHsbngNbfzylFAFP0n67GU
XYAI4xM/ckyv9Jdq0/eW1y8PpXRkdAt9m76JREXPO9g70pbunMeziLGuS81ZiWVv5QSSsyr/2yBn
73Xm8hoGIqh7TS8oU9oV5SzeQq/BYxlZDpZG4vUW52Gj90LsMVK/eaY58HSzzkGbBSa9fDcFQqEJ
Iyg4xIbewyCAqRlUyf9fB55wu9hhmjYWVakiOoU3S4Hs7sThwZ/slmG0EEN9YtbrvqqsOlRxtUVB
JCSgBrBwlO4VdyYDX1EQiCzWPmMGOohh4epjFwVPdjii61aHxt4v+OqeXNCmFiTl3z14y1p7CnfV
baXKMuDySQ5ealNjNArAj68oMB12xhU1HkUQWU7EY9H4NruGVaqJmMOYaxzTIgIwJBwtkjzqc4eu
sSbtQU4HrIRN2XpqwvN5ehdjkoNPaPh/8jn3AeGt6YG9/7BRFhBm2FqevrtgGTAlEtuLEuLP1Cmc
HbekyChnmGWBRYZv6pX4lewjgHASScM3oaBOv6IV1I+2lokgWhfE1HZtWLWyROnVRkLlbXdXgxZQ
sFUiDy0RPMa8OkNupyRTsbKsWvBh59Qz0FzPxdSpY3zh9ddtsb/JAkvzjh50FBoCE0MjVQVUVDjz
79GYLmoSlociFTH2ImUWvm2Z8NXs5/HANYWWg6BSZsbI26D8Pe+Q7BWI6rKvYu8u7o7iSqDogTgi
eszvcPuc5Jjbksjq716m/iW3Px9UURcLpJrveNGf9NW5IjhClc0rwcN0kfQWf0Oith4s2efuI1Xl
bFr9Cf8TbFiGSsed77ZFE6LFaeZec200gSD3IMZBrV2UAImVpCV5wypudR2kxwcP/616N5q+zLoG
/RIuzTLGq58oRN33CUk+FEVJcaFEhy2mFmsAwOFTKI4YGwGgd5Al2BKzIzr6p/OOMjoXmQmX+ihI
U8tQLVF60ozckeamCyPdrGxnIsFbmUiIYbsNi2J7hbHfLRU1ksBEf+2WGyfzdlV0PiYsF/dAvSyL
7rDJPmG1PsSG4jYA1gZw1EOoLD9mF3oGfnCyXbNvevbvWC2I3SmZreawZwj8W8iSUaLCyspicXL8
eGp/ZkOW4UJ5U8KDG/qAtr3fkIPJ9+rUeUZH9RdM3RLHRB8Vnv6gc/k89UM0hAJffK5LUtsZDA+h
Mc0QSQBARsaRN3Wi8H5peXZAwrqSV9iviaeHnqKZ0OMNGxSVlG5YtsJRGCQDb4GBfUiMn+Wwqsyo
CfUtrfBhjMsS90x19MhtE9anwwgPJQgp3bLyTI6GZTWaVvVQa9IqqML3N/JxBAEe+VsSgZswnRig
1+789kzdvWbkPsjEsDnTqUXpMWM8DFfQNOdahDoar2gtftfLHxjV8l39NRs5ONpZW35FhJMb8g8D
qBygwhVvzxoqjEZwHO5u4xQVfrVWsZ0EGi0fLwNIOpbI3yyttePVHvv2t1mugLiWv75dvzYQ8trH
jJQ/3FewkjuIYLChZuftKtnjA3QJ1k1PPsTkUx/kiaTPXqunYwlqfvxck6/GVllUsTvyOtPCvItC
nHCwmyTTmtyR+zeKm66rQRswuMOlgRRxMZz7cGdlbl3BD//QrhnlSoR+N9UZi4alOnqwgazI1B45
nayycqANwq5NzQVndvKmirQ62NCaBuqojevnFSTSzi608snqNDHahdFveP5iTHm0N1q8+DHGK72a
fqhdJ2yXFy6bc/HqviB+yTAC9aJOJC0RZWges2m/jZFkeGD4O328q1KK6NfqhmgeFVTyU3YrVa3O
BrEhtyslLHE769B9GnEGo6xS1YYyZKxl9FInUm64e9JuWuzZiGpt3v1Tjm2SfGWMJb/0ObDX0Jp9
B+X8gSD9NBmKY+yAnn7vZisAXlHD1bNw6D3xYY1cfgp7rIj+lZ/2J/ZdfBYkNOUAyKgj874pd3yH
eYyayMWgJnG2dZmMaNd4WAaVDFa+V31fTSqZcSynMn6MlqeXF/Mrv/yIfm60xfjuCpmGhV8mW5zZ
638pbQmN+njdfAtlGrrTWgCsrEZOaQKGWnOa/z60QGOGJL7vcpb7r/EpaCPPFBZjC7h/wx46hvRc
bdt8MCAVPYEzHA9I9gkstpOeSzdiWx3Syf794Bhi5HXG7nhRfkbNvhJwJT6xDghm9ejUibTo6zLY
8sHmvoaQNPUI+cQux3603+9kWa2YFdLvo5rT16XBpReEmwjytYxGQSdsWFp9pHQESC0b1mp6GgDF
u64Z7aiFhNemGy5TkDQFhjdaeIy9hy38SVpMwGbIXriuXXOplcOJJ1T2z39lABicSl/nO6WYe9d1
4s8Xm5QpsrxJ1JQZ3+NFHashZtUV4EDlPfd0MeAwTuwt25KAG8fwKvIjEB9aXWSCLAcsPEJpiyEh
7JMT6OB/TqSErcowpYGTlBd5e9cbrAyrra2mTgCPVMgWPvPajAxpZl47m40KAoifv8U/xCz5krJY
RU+ym78vXpfhwmPng6n/vNL1nGymbbsVokj2zpqwso8O7NvA3LnYP7l6F6vdCyVsR/epBD6wYrWQ
4CU4a5jcHdzhm9/NvxGu5khfVAh9T2S8zo+mvMFc5MmZrdr+YNm6/6eP+B5fp3Kr/lNanZicwJO+
nB8XpO7rSSIpPTfR6Gg1vIlSfBBcMpxRQyCbiTyoKs/SNdmZxy2xWCzfknOSgbJ4424re5aJ679K
fRs6330krCgpSxGhNpWHs0flw1j/vTI0v9dgs8p58HkwljYeZm1b4GUXNTo2AXa/RHaEdlMBBY2O
8bz8QMYn2h+K1H1UdVLfOC4mPzw5aM3+r0F1uL87e5Jz293FTqWDAhRHzgeGnFmItyr7opXVxcqX
rr8fO2D7pExQc7/iR+nt/JJsgIznMbUO2K2nouAIkVKC3BW4Ow/GLpt0xNdWgNNe+ai0F2Kg1tzX
N3HPzKixxDi8if7GnO1bSpbwLTQXKNQ4x6JHtKDw11XCHd7Dj0YqhNKRsmAbHcUVPCUcSrNSg5wO
68CuQOe8Dufcqx9s4xrAbN2mp1bgqvtu5hj/nqEtCjt6WuGnbuILCMoJs/T8X30sPqbPcW76u1iJ
1B9pYq16ulWliGZX6lk5z7DjnltJAiMmCEDdeMn5DAQP1WrV+XxjznlYNfWBe6OC0ueEIFmLm5/+
o9/wDhc4eSaHGX8cbQ/OoVs0yDT5YBahtihu9yAXOgp5Z+O7CxJXaNh+PM1eKXmvb+zK3e0nbzRt
uRRGDb+hQvBe9WUwpz6iU8UmKk4/xWB/va2f1K8YWcTudun0uCEhjRU3ue0pg65qmkxc0PXwhDY3
awpMYnNrKXBnCT8MFEtrbKNE1AmBZfCbADnt4EpXR2ary/q8jfDcD8kv5Z0dyvGsi3wUZhOwCQJX
kDZF8Hx2rU0895qy6YGTvGjqSD884F7EOmJM/zetG7AP0yEw9QbjIQpEiDKEfl4/kQnTWI07OoBJ
2zU2KOhJhbXVKrKZcI2P8LhgaxZCHVrTF0e8X6F2zjIAmw8/+cLBw1h3K6vln3Q8EL92ynDgrzD0
hH/JYrFlJ4ka5B7exRlIArkLLJDnaBup/Zd8Hy9QECcf7v7giLsaL0lAQHZBSyKnHjlAs0udxF/q
GUYpjZsV9nxjvcdInuomwFJWemgaGYq1IC90/tuC/iHMc07bOfmuXysGVtotMOKJP6V9EhcoV3fT
TAFVhsYDpKFvjDLeTnq73cuyZ+cZCLNq/4qEr3AoU8oAOojzLvW4wbnJBvFzBz99ZeoUgn1hOxmZ
OOvVrN0C0wMNgSqru8XDRXIgbHI/gD+3cFoU8zcyWhLOxiFR3dE5ktsQgMk+DChM6Qh5XmUBfLD4
WXzuwG5wRCQVrWcbZbVNaM0lhODpjALlweqh0OWC5/+rhkaVA0aL8SZV7MU3xvrqEPE1pugEIzer
NqFxARufzu8ZFJgX7aX66/XshSczwCkWpVzbqzHjAauUU9X2TpwAv1kpXIHrsh5aqwE9cchGec/u
QUi1keC4MD5C1/VJZLFgiVdwoCgp6FsGdAS1E/ldPtyXxbmo130wZ+T8Ldc/cF+m8yfuOSk46FOj
L/vMxqcwSFQsCgb2mAHwrv6Y9Br6h1CZaxUGXxQ1/WXxkJP7BAf3e+sCZAVXdFu4QsJTLsKHEU/V
KMbx1uzXOtPgcf+KAOIf4MbfV6QezDQqtmfSg3+OMuxDPS3hNuSsK7q8rDs7X0ptV5ujs2+Eg9A6
O5W1UzAwr1zIVi+IW6INCrODxSoH+THB2n1RjBEylndADNQ301Qz4Yb/vFOQITYtfg+3p1T+2Fo2
X99Kt1ltA/ciAayGvUFSRWFww+xgBztzdPN8zDzN9mwAB3Xw0ZiVPEMDYyE0D9Kevt4W5lTfFaZc
un8Bd0CE8MJgsORKFC5SzTbrB+SOUpHsJ3hkitomY8eXSkbQ4w+l82siQ/tViV+QfJM1SEkXYhUP
Bgnrwhstktqx2P4avobL2hlZ3c+hAi4uA9AMF7pL4r0/3HW+75yPIKBfOoEEIY/9+mAq/Mmf4gLw
iH6GyTLGDun/1heHw+pT4G0kfMI58LfdfMqQs+wJlbiGVEu3kt9gMc6xi1aHaNNR+TKEqOPQRh0n
fupTsRoDxVmEejINk7rjNeOHZrXdcfhG8M1iTehVTub4KEsJjG6K70V81hmWBF3NK52w1fP0X0I5
qgXDrO/CR+5WebNLZ/qLaeIDToVRvuP9Jyd7iK52n8U+PvieilEPYfY2HQEWxGbld/Co/ulgzmoB
2o2BXa8Qsf9GH4a/9OPlpewL9QUF88Y2vQ8joEfdPxcT/ALBG9fzrrXPCo9I4MZ52RbacT9xvpOD
dBY7BXJpo6Z5oN9+ETbbwUOlZqgKzEVzYTIwvopf/MoXQ0cumA2qqSYEwCySgkWtJhJhZybwBSLl
7zMrQdAKucuUXetqSiIr0ipD+Q4njxi0O0D7dWC50ZSPXTPwsSk1v+KnlTFr6ApY6OwPsLuLVVMI
5GLvpiCk8YvJJCnv0q+fAEmf6xVKp9ZQr6iBaLHG4wrqkMCHZQ1jm1FAQml2sHj5YJWH9m6m4MG1
T1R4IM0RfeLHwIfJw9kvjitrcUDOA7Sg1Cig5weVlqx55TqGszHAaQYqjyYqy2Pb//h4Mk4et5lE
stTwozHXOpPlBpLd1GvnikDUBBuh15K7j7+F/EXFPlZFrK2ZCOVTlEvdeftp1AVIoWx4fIxcm1Al
K0Ntc70MQ+JO7eaog4Oen776Y0gLQWDHS4QbP5W1co4MXbM4vPoKwOnvavEeF6xTwAFLzAAYcqJ+
f6nSSDjAAWM3mkWhaQFnfNmKRqMf0V7+0cl2Br3Zv8R4Gp6RIdROQEaA5dcfDBOWcfKG6CthwSI6
jy4yG9xQYQBwscFmpaGLrfsGnIxjS6tEZPn55pgTgrKZDfgXiEOljfSjX4ajxLWoePTZ/sGZGXF7
Od0pY4YAidKGWvBEOKe0fXXvf2EUOZLf+8ERTThKJK/gGS3Fs3FEuLlh4JARkykRwtYaJasX6hb4
RJQit0b0AFebCiVxqsXw1LSZR1H1zKJKp3SB0ZKPN8A/DFp/oFznyduCVfy5WXmO0oQfxc1wz58X
V2JJGZaooe9bogxqkn65tbA7uD2epJMNM189+5u3RIwPSGATdOZt/oq15SHl2AZDCFFH3DcbeY2e
I59pUX3rxLP6AV0TyBFYJHOrPxAWmzjStPWRRz+90Vp121mCO4NEODne6XyH2xGImW3s2xAyLX89
dOqSspvrfwMZ3uWUztOnyHjtExud7wxI9Q/HLT566PlJ5859PYc4Y0eEWWO5Cm/BjYa8sQ7w7xfa
DtCGDEgWh5MG0PEncTGeud80aWkogHnQ+5lw1HQwQOWuJU8TdDmZNkbUjSd4hFNafH7RgoCOpHg3
i6Uibl9QDLrXPZ+BbdGiWb6lc/pUXX7rdbA75ixf59/Aw1PRHgNIs4dRWjK5qLsvi44s01TB1XdF
tI/jYIfuFgTovD7YxZkQCu1HDNo7fUiVd4YgvdZp3sQ+5z84tGgt1TZxob3vCE6pk7qzmaf+6FJr
LEn5x+tI96hpDGKVlTi5LVOAwZj6gq10ouBehkwhfV7G+bhmb4nPbpu+zrE8KYeKhSF3WrwOeNPI
rlSlHMue7XS83oV7a3NvAxAkwhIkGett7YuXnnBX4ty0JVRfOdQrIkY+Gvt8oGD+ikko1VqnLG80
M8moCoQG17W4PIII1tRk/aephgn4/965Ns3nUnp59pzjeMQUO44jv7oUddLaz5ho8y8aVn+PgRLS
WS6cf8/KSdlrGoU2umtviWhp4/huajoXq2IlSGDFci8fFnwO43iR3euXscPJ7CgT8DlC8+2M/xt7
xrkqOjdq9c76Gux0igwx8K1ade9qHhM/EcX+sWVTWTnTcbzSB9WfcI2c/jOT2pChkTGi41Plz8IH
xGsNvirTvV0eVkknZGgT/7L5QVfFavZ442bedV2MQlhg2OoDm6yCJouCjAqf+3qDz1chpAb303GI
Mg7nLZGlNjDptkD64zjkDjrEgDOEpN6UsTb4t05/0b3nhDyOPokuW/05YXt0qoUuVesWka1SWwul
JvXi4MRFrJJY/Wjb6NtZYWlvqIQFPAQuAylfYywWIdQ3GVoJn+Spr/S4y5t8DIfCHETQyfHAqfhK
q21Js4P/ya9EZRuK1RB/w9/Cqdn3QEPGJc2bzeKHYsKitariPXuNScv7aBc9zV5GF5btuiM0U0gp
r4twtjYzkLBVPzvWWu6xcyKbaTgyRfc7U/oGF2byioYWOAfGGxRByteK28Eo0k7L+I/C0dqQwovj
t/Fi45zFgyIWKD/Hhil+h1SsKPjI1Y2Szw6hluymkt6V5kAUksgMjmlRMSueFmtySk1Aa1WjWH24
1UR7Fd5fb+l18ZApSeEgxMQq1/z4muemUNCIs/MAxhsW/7Msf23K6mtNNwXHVTMtxCVh1hAuEThy
yfigQ03pNlYlEaAOX4C2O/vIKy0t0u5LoIsfDTSoGn1jAVvY/UUXGBosaykhg+ROJu+dpWvsAhEL
7SrdOIBIUcirXMSGmZAcFkV14zu5bDZH6eLfE6s3GSRfZeTFxwQVjcDrZDTWB/2A1jQfPs+O4ttf
VKANeBhJEp3lhiLkQtWKstAdVrOmcoIcKjCixKv0xyZd4+qYaDn1PCUv6//Zt0ze6cP3FGuOqWaj
xiW+emj8xU9hiaT3d6PjBgEprjKYlXjREH8JYfCo+54LIV6itqAcPbJ4mHQI3Mxst9+sLqK3nxsf
VVFd8CfDeUQE51ygmtAGtk+rUMUQiA3JrWfG4kEKBn7hc/E8kSS6eLSHM+x/NpsE//c7zZ2YAp0t
tGFPoq9hD9h6ELx4hxGp+S0a9aW6F/VyYu7TLC6kw6w0nR8jEmAonFKxRxH0hC1cXkaBhRb85Apv
VfBhdR07tX1WsmL+k4k9cYfRjSSKrvT/Cl1Ls6+wj6EmVbDyQa3C8k6O4F8q0kqsFTYaxGFjJ1LF
iIpmcQVHEoonpP3MG9rrQ5k6mppusOUSbEaoe/inwTFKKYaq+OHCpMAVrZkwmWcVcTObNX+so3Pt
jJUGX5fKbxyx7xpqE0vrrjAMHilD1Xt+pWJzy1Bg3WgdUczhKXszUG5tzox1Z01q+jNapLVggTUI
PQIQc0wpWCI/x0ikHUE/03SCkJID6Md/QMS4ayd3WotmLyA/E5a8XJImb1jFaYRLIXvLwnknciGg
QetqZyL1v3fp6NnvSApJcEpvGa98mBokgV+fjm0WFrqXwxHCrmJh0U/MoQXGLZTYHBGLJasdaq1p
SnsrN9hYmw3ZHP2WFR/Q9ve9G6ZAeUu8rS7k1gpx2tDShY3v73DKrU5Nc6thp9XTZq0U+X8YDwMj
E2UIcAIvb47pFj946Q0gicCfewPZoWQSR6vm6ifAZGG34VAQ2KMWBekgts/2BFWgmaBkCB0Jppwd
PUyW5ZRQ1COkuky66UK/qov7TUr4YRCdSQvzNuqoPjQkJKrBWGJYoN/hHoj+YJVUXdPPFo3BQMUG
Tl4oqtOgVzcEvW9M6nuMOhlUiR6Yzv0caWc0QSEdO8WqXrAh0UmfFQlTgLDEY6PBBj/pTAvCjOYX
N+Nm//7hhfnKX9JafcOrQw8aW23hDeKhMeypfZBDzQ5jwhD+dqUwuqS6S6RugnUW0dvZthtomoZo
v8ZCz2dzy74F0gZeZNFELn6VM6NhW9HVxXWYP/8JweHI4g4vuuPNzljgJIdmeqh+dvAWI6CBDRl6
qGKnKcrTiJNMbo5TzrWt8FjVlDgzMGzQljgikGm0yLYBTvvTDzuLrAcvLmAAi+LwylfaNGAmJsBr
2Ku+G6eArEZ+FxzuvK0E22YN/xKRSwCK9SQ07n7eKd14a2Qrk9+/THhWeY6VKuebK4E1Ekt6wvll
NBiHyDYTOuZipHqJDziIjJ9McnobwZDzP8p73PUXWvr+vh2gGu6G2wjhNcW31UHUXIDL8MoeGbN8
GfNNXbckigj1ytwoDRvK9IscTvv/whxTXqSpm6ZEC5N0x31vSihizwjJWfBx0zrbE5QxljxXgMa4
CWlp2lJoZRo0neBy0SxlVrno5TsnOl9jnpYoCyTGzYKh3dBNL9yxjJZwyPcwYTUvl1S5I1xiiO7i
EEOT3uCFwL0Ygocr2Mj9GaYwIM9hS1yk3zVN/0zEVGR9/uSq6lvuc5EhoTsEeLhS1UmUK22xtVO4
guoDD+8qsjGzqLk/bQMX6X7iuwbUVvnIAk6w8ECJG2rumhBXx1bn0bBNqR2PUpZIMjYw6mE5R7I9
E1X5CiPP+3svuVxuhZC2RdzMYqW2cRcU9euAL56rGVb2E0nBLF6G4NXcMJTzPnp/63L532IlGgZi
k5dpy1tjlPrk2wpmRfPuSpSPoJcEr4VGtHAVK7AA+Dw1M63OaPdEoVwrhKOeykV2fFFIgzfgtf1v
JAbzfku7aiDhhR71tlCRWron8mEkO1QHPkDk+s0nQDWC6hwS+8+0Uk5AYDcgkTozgH/moEeubT4t
8bYCT43qBuI+C7Q7Vmr5eMu09ZmuCX1XIQXY+FsZjQIzmllnwXZvhPu/yoliBZ5za2sgmggCfxbK
uXUv+0nlpmj3N9ZFwqPlNqMFLaWP2y/tE97srqox5WysjOWNJ/wvS7UqP3fF2QJbfCJYEmBBKq7U
Omhdago9aPSaF0jUln+FsXZuE20d8Y+pqkukH5Os8N5UoZMp7KAxkhCP0cEHERf72njyH2Vqc3gJ
4FGqau9n1D2oR43sEk35+OZmSAq+RUUguwZw5UleKfFLln8p/7G8KYwHqdBj+9zHFIbfnD63tYuY
M6RkcxV2TT6PI0jbOCvj1Lu4+ZUHRSn6TrywEpz6acfmZ8Jqpc1pPcCZoGPEatnGuIXH/7T2q510
OG/xUZgTtHRqAhifC/RJmPwbnZiAYhiILHqBcyZOjKpZ76feNB6A2E4Ig87fTWuWK/NCw7S9LLOw
JYyP12tXCE9HS6rBH535IDfdvAIaR7TcrtUsnFFuAdsHJRzh8PakmvPtD5wysZbgqsop3Kj2Pq02
uyipnQue9EKXYzC9twYF9WHPuOWeoTwvB6rrIJUWU7g6zw7+DiBVSCok6j80k4xn9s9xXML2TMjK
qp7SqCZz06rjasTxpLZzRiIY26ZVZv+E+CCuxR/97xS8Yka0epe5OZAxV+4gOd5eGncM8X/0KwZD
6DCWcfu27oeuE/Rr272q5rH4rW4P8UfCDtbRydf0oBuw4w+JRzzwFL0pe9/cKUO5mVSMFPsD9j+7
muT+u9yijnT02LRvSbJymUSowbtMvJjzwVtnf531JcGAHPoX+VpFLGHSLikfxWAvR3rgr1bm7FdW
UjrD1znvJ4Y6EardMtKI4U0bEt6YyusX8K37U5YnqQ5Pnoylr4V6GYybu9PnMGsq8woDvytkU6Zl
8JrP6la+ADIzG214vd6myxeYreO+cwm9/sKQ4KFJ/OhYD7Tz1qP8yEu/Uncva3CIUJEax6AZNDkJ
ZMFanii35fhqcJzLKLFFAbosCgmGtrNMotRuQZM+1ZypUo2YsxynBbqh386bHHm5ZVBDONkpP2kg
CxUisZf2Tp8uIcP/UBdS4k9yslu10E2kyuSLsa5AoH4UpBfx7QSiQMmhh4088SzCpsBBjIjRh8zQ
d+oL72DJBA638gDJ6AeWWnYbUINvWKWk7M1L0D8GEznm7EVqY9ZDO/qsZP5FKXpAqZ19rUw5boOE
QPl2y7c385L3dsBxLRp8F3fVajMM6d7HOPzVgak5uVawMgtehtYZuSO7oJCo/NChmKosY5/RTYYg
Qod2kEB47bZiggAjbAxhbEjShwsGEGUxJ/Hah031Riot4ExtZMIOSxqbjEpUVPQRPiCRFY5NtSmI
evutdCupsPGOSu9SBuN9nVKU24BIjwrJDfEo7bHHXT1WFvFQAwrgT7GIJ5/TCRBU7CnfgrLtnr1n
L5lCzXuejXjltPFhAaJsmWylPzHUB20aJf1lWlq2dHH0c1IX005kDcjpXDtueeP07F1hcBNz6juS
GoRD7Y4IV2LdFsTJjbotq8OLnY5gyoi9qapIGUunCUAiHPewPJ7Pcd/3TLDdUV/K9ulcYcqQfz4S
cRLfiUN6eJ0Py12c0PKu+QoAfTD1oQLerE7s/Yu8J0oGvhMoL2iGkJKlaKrcAC5wjLh7vfqmB7Sx
LxDp7k/XX11XF8c0DDuSBPxa8fpPd40b1wYG3U7E6Oj7FF56n0nUg7G2Z3sNhayFOr/OUM7jPcvl
imEvNLvE6DwlA7oDozhe4DwHyBhnDCNOWbBu8AKBt37KYVoJj3syb7qu0xXSxz3b79tim3957YDQ
+VRIYsfNynhEpOpRxX3ZLGTJyt4EJVbVfsyWjOdNUs0I6qQR95y3E3Q2hNpamutcwsryz5fcEVk8
ZOIliZgj4KnOYSi3EL3MKQxt0dPhcjL7bSiSFyCpg5Sfogxi9SMhEojr8KtXSgidhl7fzhS2k9w9
kSKQZRoycofpzJBk7lvWmxPppaB4U+mxJnYiGsBuxAY7bdF8akPG6tmtVM/nSH1euBpQLeaJCasp
WaUKt/93G5FjaXn6D+E3K/8Nzf2/n9UPqTtO2edoBFwvL/tqTQH7B/ZC0mQ30L3SHkAGzOlAKX6h
1cAgf8TkjjGFJaNnMPfSMhYH7R7CtaxTbuKLsWknKXrTe11aUQBM9uu3bbzdIAAzmJ4eu7qStVLh
D/TUQBgUNIJTPxwQMPvD5RWU2HF2P1WLDCiHGSFq4DFUpc1J/1Xbk1+XJtfXa5g2Y8qiSKOhcpJC
gEtqsNW55WXkyRgMX3ojjghnkNf5aSc1yOV051tQ4UHytTfwznZ0Lb2P7hKMUlQTLHjLniU4UY5V
oxfsYVNYlNx9UltcRw5SIKyJLaHkbktMofdtSbp/rz95a5cWk2ANN/VT5118HmU/y3ov1yjWIODX
F8DCJgqfnGNRSiBWhaEK5hVXULJ401ZMD6rLbzDBJyOTf5hTlYg3BNLxIQhst0D1AjQr9JHrK3eB
CiLms/Vm9/5eMOqQ7VRcD9Av13zaem+fwUBEmDwrfjHrfbREh2blOU0atrrqXZ1OiTeY0UjaT4sd
If1xH0XjIKqReyhFjdBROpO5gF1azvlCerhEH5+7nEcIeLlb+/AFgmeR1y4BULHRT0kJfobzDWWJ
x4X0F00R3HUri3B1cKYb8OI2C5wbWc/ET011NNLrZRKdelu1+FKcZKKcvXFtFjxP7UVV3ZT9lkKC
19H7g/wvp+GBuHf2CBLawSzIKcfsgeXMjF5UIdv02YFwmoHB3go5N3TEY/9MkfekZ8XxtrMfau0V
L+HmbR23/K9A40v0rgcDesy+cThF97jz8Y31Vn/Dj0jAMeAq5+g7OJQqtD+yZY2RUCEunKbZM8AM
S83Hdd+Ij+GuxJZj/bqbX9uf/mauIhTsKN0TduIH4/Hbewyaea87aLIlGznseJeRdvzZXfR8krHY
YwYhWic8Xn+msCGzW18d6oNcoLiY0HmtKPgKP13YCW1mIxjm4G4La55//6YMBSAkWwuxt1ZZMFhJ
b5ZmVbMEoTKMy6Jodb1QdJ24m8qAT4dAmkEbURxoqcl+gxDP1ckfPxfM0AKBcrD+Yjb7CTvnbSP5
RfQQYYax7uvI36d43Q9M4ZinAwPqiFueyDAOIjIA7vMq9XWJTbjYRZIjPrakWLZQ1JtB2R0/on9z
LofrdGX4peR+q+lEnqrgnA+2crFsasJGWI6uVSkRkRGiHuI80sq5jTRKn4fdq/CikMZkMBjjbgHu
w7GCgQ0snQcwYxBAEgrSKWrvmxZgYYumT1Zmf/iWGfSdGNi1umN3y2fjH128tvgSzhFA58E1jZLV
V384lEFjz8o6cvmbLgJW4xYMirX3lnvO0KysG2/5XzwQPHg41ZG2FLgyrE/Ss66JpoNsdiRdbMcd
b/fmhIvZpmZorMfdFKLRub51WsrggPMkqBjnOpeEpACZx1rn79Q7UF5my9t/Vwqj/5Wl3SjO0gV2
JOMJvVGwbZsVo++6rF3i8W1xrmfYyHhnwfgIRsatFNEZ8OUpk7i5VvLcuOxXMvzKJrS2APgb5DYz
EG7CFiukY7uHC/zWAxRAM9qvYTR3vZrGCEp5Scae+VPOzJ2kMF/XhNjDkSActdqngXQfPRk19XXS
uqSQNmOwWpA8AQzN5hzVqqDhgWbdyXPWihRPPHESMMqHIPVefMUE4uvIv2RhRQQ7N5CmQB+wzlWo
oSwpIcQAHvkzK5gThyKP1VLxbe5FTjc7aHYNZwyBLBlTrtR4dRUlzDPRDBrRRQSCno83u/EGWHCT
lq+TdGBGZC5qrBKssYDYLCMt5DU5sUzrk2Ni4Ct1BFM6mi7gmIwvQqgLGtxuVBRvyUBAwmLYNF5o
byiuL8ZjeVvXfBLfKgm4lvva7k7lnC3vPiYkDkEDDbKcsvgzb10R6fpsXLy0k6VCPaCdqJ5VrO3v
F0+8ZbK1KiRF1/N3hFXvVYitL/0LMhveEVj3MkBmKnka9TiyN7w13QzSauDJvo/3wtA0/Axyg8WB
lANCqgcRLkTjLLfzslnQ6gellNdprN2EQq+RiJaE9MXemJJtG7pzeqyGJpVS3QX2Wp2b65XAxMz8
ScErjoujX1X92ESMfegbAolUuDjNcBxuJnrg8xbxdTMkGuVTWKGvOYqqU8MhzEoWKeNeZ5zaTbAH
DEYVSK7e0k4tVKirYR4G7/O1ly7TUc6Nvucg3zI0ATHfC6JHPXhMZhKLYskNnfw6Px3zy0WJXWcU
VglaSdRYzHWnW3yVtiI5hLNEoLwWdyIvkh56PvY7wNYgVwVRK5nMyY+H1v73blp2wi0m5iX/+BA2
L9ScAwWzKqtAerm2SO7zbSDbXy7bc5WtnkKS3SIfc2HLWh5jKuafV03pSo9pydVyr5p5lhoB7T3/
qva4O4lhJ/gUmrKfpA8nxYXQ4G3O+1QbIIIB+5pJnqh00E0123kpfperaXZwKomZfgIpuY6AzUo0
dr0TvaNiPpQMnQOkWTzjNflZF44s2iEMV9uiTwr17PZT5bGAO7s7OWmaK435+kXnAeSRtNnfsUIr
adZAzKrjoO9XTkmdrfY1CNJ4wKIQtZE/MfA5Y2kPo0iuWorVxu/dprhkkRETwvRabim68CuQCOEV
UupgTDc+RHJt6UJQUH2qRpMHs0iEonswZIP1tfv+zCACyXOs0Pl7513f7jGVLlgdGRQxITc5G4fu
DjX+yyBTcY0LADUUSNkBlblarDG+AiuK43QiFScceM1JH2UX5aCo0tLouPsIESFzB1PfQ85EXo3u
eHWyr0List1lu62FBUSDBOsU+BaBOe2U3nigfAtDS4rM6ziJv+2vYGRS40F8xTXd4unnSRN4a3LV
XDAndIF/k49wRP3RZMkvUse9+3RJlUbJ4a7fcF/UO520fcKjRBRkK+GVSZd0Wh8VQNmPE/3uADkh
sI6ir/tICduOHXaywLJME4I1Yq1RPSAfpu1yQlLBNPnLMrvT5ODiiH//rOVhrUNQBn+grdiHdCZ+
lTI/JtjvTq7uaeH2iQ7WxB0gA5dPT0QcRJIciFqg+Y0GE513/SdS+Buok+sEXezC2Kv9JHDXq/AT
SZFt6hXzHjOE2eDKRH7dZfpTA3LUSyE9zNm8aZnVvMxuM9p//D0c/xDw5UgHrALJDzc8zw4J238X
2J8uMKjnuYZ2jh2ueAWKtvWru7ON5Y+AQraixh7fe7WUU5hPgQpzDO7BEjOqR9pvj9DjuM8oeYkG
L92TwJW9Fwk7jC3FXNgY+Abua8NK1t1weZ8p6KWOxtramK1Nzx1gzpV7Jf/t6KvJNsQuIqpZCloS
6VgxC6Uq/6rZbIer9bavgf7Gbh84xkd4tvvVrGwW+i/RmzUhpBQ9ofjv8EgpXj9hCHT6fli3BCGg
0LrPJ5Vtbnv+E9PLxArF8JMeMtNhsdmkHIYIlz+ibFbIvMdWbTwiPfiaMxol0mDQ2gWo5OLMUVOR
4BAiu50tCqzLYsqOgTqX2k/eg1a8vuHdZHhPVgrxH7+dVujSGnIyS1AGv0GVzegNseSdfR0INWxj
RsZ72b4kGJ08t54JuFNj4Jq7DXxFQJwlOMT24gi/bP+iqfYfgoAHuvmA9GZCLMSedGfS3Gcsj+4q
kdWB6TjIEy6KuJhUppUk/0+Tc+W4ssqUGjN5HJjhhsVJ/94qiF+9+9G/+X2TeTTGuS58/yTlmfZA
gXMR8h3KIKRbPdYAvmXEW5FDKedoMK/T1PPWzZ2U6A0MJQJ8I5FpaVnFrgKN/r6mlf83BqUvcTzx
pqc1g4mG/zCzuMpGCbXsNFfCFdb5TxckjySxEB124KDOihdoorCw2JNOkBtYb/xAVWh/J/YfB4Z4
NA0tKJUoIos/hFoe57M7NVUqiuowxtuK5cGaWxnKmdbn65mC0Oi77R2+LDZSvd0D+1aYnff1IslM
4vuXxSuXK238GLk0PBYeQ1QjAFZYdIhSQ2RI+sI3jF85VLpCbJ9Z7ts6l24h3NMjt5A7W3PDzTN2
laURgSxSYQZqY8kGN2QtV9YlZsI/u7tDwciGmv8523qm+s5z10Xzec8ym50Mh51+iHKPFc9trlXN
+vKNqp7PoKM8NBe54y2CM9HY/jBYA/8RnCrmFr3PD13FA4pYcaAhe6ERanmNqioCJw+liNdFenrq
gktS4T7toJ9z4rl57R9CTfZMo+Yi3XFoGohh3qltshzGNOqAIidU29jS6KEJWx10PGdtDw+EUYcw
Fe9k9bIEq/yg2dXkmjr/+I2TeCGY4VyDiI0kCPvWvqwzw5pAleSVeoU/Ad5E72L3Ol59JrX8ZJrN
ryLVZcYt4KYNwuFPeS+2fkLMkLc89vh/lCWptjYkFhxA4tE0d/ZElaGhzGJTrMM+Kouw2w0jSTtD
D83e1KP1IJtvJFrnXNDI4D3WleMF4XfOB09XYedJVLTMtlZ9OKwei2b+UWWvj94kbJB/4NTLABk2
iPU+pKWwQapwOBgt6J/AtU0liFRspfqxWQbRFwdUG5gR265qN51wOdxqRFFwC976KV9Sem2uHehi
bnyvGRe67bDs8kLWCHRVp7pknMphjE8WK2Abmxa3qD37DE0yRtOyTtNBRiV3qvvX5RfbHyjGyhZn
wkCe/L7T8hrGf2KTT/Nz4S5GDE00uxUszLAUeGl73ln3tXzRXYI8U4u+G6D3QRSsxv6eJZZOqmey
esYwK2b2TBCTifobeYYHHkhsnSmZUuPf8YkfTlsx6NoDMJMNj7mUSlpAtt02Ts8XDsM0o++Jy5Gc
oejEEf8Spyk81krYQFV5Wf+scrRsaupDFbfO3EPzqZ55Ne4W4KNDMjULjEjYTb8bLtzP1kDNlN+f
7/DbdrBsDJfewLGT7L1OfbnHEZjT5QhacgzEwmvVAwdGiw1ZUCi8u/5wzQCwN2tMjAJhUh2yNLzi
94ld6wlNkIGnG+s+IFhxbkNgE/nIvSabOu59ddRArpv1mw9Y+K5WuSVzQQJ02DF8tv2j95+CzP/c
H0Y0zGdB1Rfo4qQGEc92ctFfw6os+4kDbmNmlBfBNrBVcgJGfU+4866kGhIb/h2QcFpsyyi+Knjk
BFAw8GIzyalEyC9qRxNzOp/EycVb2degBgPDvZFZcM6maEfTcVc8oy60jjkoSfW/Izq0heZBt9q5
BKchbqfjMNde0vloNLyM6KRGZ0lvHAyOt6GxMadoRWaHZATRvy6bH8A4c4mrfck7/Wj/kiV4S6KH
656A38NDsO9qUDPpvPn8h7PFpeg9IAO8CS8Ic4X6zwZ5l5qwjv2m2Ah42dFzcOZyAcOmfH5AZ6kN
n+KRphDzxYMA85+dW4MDCcpuTlHyJLGH2f60SMYs9exE9sWyXT/X+KmX+eUWycfHw4y2eYZF3nzi
N+b4B5sfsi7ZBvRN0UXmPXwVXLWtHIo89dchSThOxytT3F2tPOhk/Qwd+tdqZzLWWA1Qltsisvmx
ghQHyMGy9PWORuSddzKCGuoyGoZORTOntZ0RpIVdofyVC+TCFLIZ41v8PbBqcoAMK/i31e3lm/ay
q4O6kZqcYRga9T87C1hYkmB+JeK3//o2EMTWEPRNrxuxtlmAARJ8PB4V8haPM45YXx+2bPDoNHx7
ySVXLRrRABNcncbkKxibZRxztyT0MaamcP9Vt+tAIVoVOphw6/W/zWwyJJ7ymoiQKuZeKzx/5xkq
+UUVuF/SNbA2247N0AYV1Kq2rILkcJzS2wDXxzA15pCly2dQm7TnbNl4h6LBAxa6Y9HHiGRyptJ2
j0HJdBTpDOCgk+Nhezqc9gjUTjIky+Bb+HDdBVzeE6lqEhJV53Z/a+lEAQEeJNXUzl6CO8qIsXci
6twjSA+SpMeU9aMDlC7/3UYqJV+0DSxOK4CfAtPP3ANNQ2IUzTzUKd2HH7h35VgGEfBNM0XpL3x/
TKzOYmjXMh5HgmwOu6V6OEMNXDIsDQbR6vcccMzI9qCDDNPdcG43xPUyM42Dh6+lYac+5xD+37FP
zvdUmB2S9aWtgcKwv94wf/V0VlVpQh3MgdoCyBR1JH1k+hTUEUzI+bLfEA0K1LDBu+FsTmX4y+q5
iOOz5Hcn9JbquDwjsf7jj1T3+RWAy1kfMphxOGKxVMrMuU+RPw8pcHD0NxZSvZ5BNmG+cu3/uBty
h+f+GuqmpCbGzJGtcRa3caXeuWHE3hS/dM2ziGlEHLcGSoZCQ8wmbjrC6RsjTwjLBDzwED0bqYZ8
NN9WwITEfqAcY3z2NIU+PjXDIfIyfBJkmHls0k/G69Tt8IEuRacHUpqRcYgAQ5iHw8vUGMmgGU3j
cmg7CNrudLUaC6IOlmRXgmR/Woz6m5OsN/Pts8DkkoILdcDF0tP8FVvtesW1OEr/N+xmX+SQObcp
S86byNHXBHeuBVmP0AvUlanFXRK3s2IjIY/QX0s0A+TjaYqsJXf53dARqj2nywNdY+lHCUDegZ+D
oeGpn5AKgqCHkAEGPt4lIli16fncRn53Ch40ryIESZKgtRWk5ebnci3nQMctNu+VyiKTGNM907Vl
QQIoNuMsJBz5nwADj7kfEnisem7CqOe3BLpUlLsOV9OfW9kzwP/y31fvsxigzwtzBYj0Akr6y8FG
EaGdTcGAIxPmZzAWd7Ly8ztIzhRzwkbCEPZnuWTZmhrVdfoxXxdE0q54LLreitqSfFxo+lNw4cNG
8pbAiBdA6Fm4Ygg1RjvFMUn5HjjC56Ble4jvYet5gfEpKMD4c53nnHzwaKl0pEfhwPT3nLSezWRo
SVTombCbGyFVeUBY9++TGkxQjiT31w6iAo02lPvuw/GLAtGUb3qM4vOjzzjJHF5E/Hr32RzbjZMP
YTgNrCpHuFpR64/d4fdM5WyAieMfxYOFk1kUYg8MDA7Ywg/X2EqwNS5CFcCpfUO0joAhRHou4VH8
A3pc9nVPLk5pWwaVVW4OL765/Ie/U4cB+PTUKPzl+iPgdvliPwFzq+OPK0DlKMm7YgLdU+BqyQZ1
V28dWX8xCe0Xrz2qOT1hvUeR5NdeJlUxrrv18hFaHFqM1sAtpN0kk3HuVRxEl0YvFNomjBrcmcI2
zcgt9CEujwog0zg95JxS40h87m2IIPDRwqh4fsKgxHXpLh9z9W7fdjTTQyq9RgENimxSDUbjXoBV
7h522ieNXIIDeb182g4KOWr71YGjGhmFmFi/3ScfndsBoCnya7ZxwkEzr7O6s+mVolNmTQKiSpbw
FSr7nrJTJFTHn5i/Jv5+ZLSAl2/ddiloz0HUm9DlUuJUw52bYyOGVStBaDLu0by/cEm2CR99fqtz
vui1+4EJdr2b52IEFiNi4NrF3u/ORYFaeHDHSB/Mx32MAEEUfdGwAlefmwxA7h/QChI0vqj6ViJ/
6mH8nERZha6NxGuR1W76apcJaKY6ZD/RxfcqHI5o67dmzIc4uoSBU6cOl3pXJuni3uKQl8MpGXEa
PhVGGb5n1Si3KdTKsCckJV3pZ1xu+RS20m256wg9DP2AFtuGxJ/z5rufmi9y1Lptwk2ccPhdW1aF
Gg3YDf5SOMiWhfZKuAmmbQNXTO+LpvYbVovyT4yIDfmumpegKrBrYz6Yk7Yx0vuppqoTF6Yop4XK
3EUUX3CROWdUxSzfP3korg7Th44/iqNWm+6drVPsv8bsYYDWXPxK3g/IsNubaNVFHAVxz5M+yR+G
NC5xnx9VAMMDsjmIXef7/nVemq4Lgj1Ayu7yxMJ/PquoBQPyx5A78x3pscZEAvMQzWsKAVWVfC2c
8AojDf6oM5kWvwTV0bGJWbx7mX9ba0eGN0/V/WSPqRRHd8fjT8fHs1SPUWQRnpZpUjg+APO1c6/A
yPZcoQ8N6IisOyLZ1f57VjzEg9vgovyfdU36YcRLCetiZiFjJun5YA9320UMJI7OOCfnKHray52/
NdhZFqn9vMN4m7S8rrWEiqKoURLw/dzB4Lrzm1iRtGDPAOjdkPcepvqL1QhYTbt3nX62DkGcEKRY
tpjejfqlIFcYshMor06C2mrnz3lyfrSMWNv25Wm6sivOafOGhh70uoOBALv1u34V6R80e+bahPC9
FjUBsKN7aUxxqgM5de9xA4E96V1JiYy/n3ljntBgfATep2p1cUlmBfRC+HqGCitTG0M/MTKbIvCl
B1E6ReCbscTieEOlEkLdnh1urXF2E5Z+k110lW9QaQFYaCpYL8RDPq9LgTmRDYx4XZ2aqWQNaLyS
3TAyecL1Cd9wqqCGZCz/ApsFpvibQawkuTmC+qrmEQG05IXj0Inzw5fVYN+//5K0l2TA25DkNFoR
UzRNnY4pHzohkObpM74C0J9DJEOsg+Eq8HEvoeYZ52YSTIbOBhAaxlURjdRPVrQ3NfAYPbPkUpYy
6/xnbFmQ5yS1DyCCo3+w1tX86/T4TXE+cN9aZvM/vh+X90u4DkTCm79gDz0grLNdUIgv+cGb1Tbg
kI9+UhGYRQJYCaZdyXVgAhHyiESI3Wk+T5YFZSoaFwCOufH889YINP4inPD/lc0rpJgTfzsTXFEU
1dG6LUxlDL2Dr4aPYHCA4Fq8XgE/W8iKEX7Mmje5DW1eYQWCdongo3YgnVQnlYzISH1iETBPADlZ
QOm8iImshkZFbEY6wKMeVObKOY7hSh9c+6ahyJ/mGY2XFlAlPrJIuzeGaKA33SRP8/hhOYL/Sflh
LPTsZX8xnp17UZkSjqr+zZGUnT3DwhWF5lAYAQsR0ywlkznI2+2IdbPSD6tCtgtL1qASiLoyA+H6
R+N+gG9ZIfY9lPjdYYOGWKloIywZ7zdRebaY3hJC6tc/3dR7p/Q1Kaz7o4aQwrUrOXTtBWETl2+e
HajyOymcf2m+5MxJhjr+aJkZiT09FOLoKP7+DoB7tIfNuTAgC32rkmYe1xCBc3wVsaFr4SYLuroF
JiP+jXKpDWP4n/BeNupAMNqAUuO33WiJ1G/yv2I8OaeqpE4kUq2qUKNvJ9tXuy/2W9i5Q+/PsSzN
JyHxHkO9KQRWfW8QuE2vpBQQgIjRTlt3V1qWCHVZrkezlFPd7pAsswn6AJBNrFMZqgV7Y7FwUZ/t
qR6cwRBCQen5hSpZjFlv0Ab8KM+4xcpo4YM3jo+AWyLraobsfanZBckdIFAH4BZJ6aCkwUqioG2e
YvoICaljkud2sgNUn3XcUd7TSzSJFhQAeBRG/UuhdtK6HHc/Wtekb44awp7ZI5o4exS0TuwZV2rX
RX7l5YEFFBSyBpJ23T1+sRZKYcc9fQwgIssafyvKKN8/SnWCRGpAQOQb0TOrTC0QFdLj5XyCeOju
fI8QlGEWcFSKsfd8YpEiOiTWhz8phTBLUfysktr7WFvMfIHv70faV680iqA9pdEqDy4x+t+KEOYx
erwx3ir2NfVn0l3lofQ1QFaEqmo4DCGRDERT0ZIrlWrvQCkyJ5BpsarcZmCfrml9tAz2rK05cqev
YpNQseiMkqRSm0raA3F7oW7jfQSE2ohfGbKnRm0OL2QtPEl84IyPa/SZSu2H5+90ioiAtMs0gnIF
Clfzi56X79jSHX5bPjdl5o6BdLBuqCNxpr9nVh2KvdqF0iarauZ+xvMNYacvtR/XYtIe+mWaKOrR
fMC0L1F9PVkPUPDrh0crTUFAMro0AKXKV1ylhFx+UymkbjNOpI/SMz30AoQIncpeCJWuc6OD6Ecl
s1Ym+I24xdKJb2zmqEu5njHOnMtnF2Cs0NvcAOqTddU7DfQe2uj77DXWARE7NOU6kIq1inYpzHpO
v5+ONDjW4ZrJlf7OkVXIkGXbYliG/peryFusm4lYtYajgJrLkIps4Rg6tgaH/6HwkbcZbVx8TQ46
IpYxHTPhV1LAx5meWMfGP4lR3zg6iUea4XIHoFQn8LzHlyhVZZ8ilVM7rR9rym8/T6FBr3nVIfSX
wVPvpx35UyfUdSLR1HNBZ5jRLPfh45hXYmvxwv0F/4U7ok6ytVyq2BbN4B4KIIJ2A1ek4i8woSKs
djzUsJjTTjpc0tGCDNpF0a+5+G/f2Lk/gPa4xoNANsckhsjthc2H5myMERjGxwlxqR2l0G3J1513
N5CIxDlMZl1C7WBzVmwHUE/R2cAlf9k4p/0uRTfbLw7bLAsEgolR/pgaVmCOMcryzLNBbytCdvhz
q5kRqkl1/PjTikZQ3TKuIE8VevnXZ7H2JVZn0x24zlgJICYWI4W62IbtMqupUsh6WhyLnAAS2HGO
3PpZtUOjOFspU0UnwHBoXZJNmCJ+3d/9iiaFK+uk0+3/iczPcOyWyUyTsqflmCeVOq42EgRtYKo3
3Zwpx1yl6Q6OCr954r6UTBapbwdanpzT4etZsWPFmOO0Cxhv6bcgUqX8vicMzlEU1rtCFOCQkKXN
WXPSvSvM5PiTlCZaHE0b59vhwUnxZwUTOzuZw2Au3Fqk53cBHUmAXFo+AKyhUC7vezCdZMU1ZRe/
P0JA0G/Mq2fAYNjyfbVMgzfFRGZXicavRJt4NYIgXYBMJ6C3SnPr+gB3MzL2lEfhzxzfTCBlvfNg
KMc9WGVxrN1Uhk28bH4/Njip01rYxd6zn/yXHM8Rzi5wGIg5C6OISG1TlBgl607V815YSjAU/G+T
/+4FfGZtHuU2nUC/ThE0+WvisKaA0cvZzT7VxYy1gZxoSzq1097biCaeTF+Ssref1aXlKUrvmid3
b2vYPsXPoUgbIFlqa4836MCunHw+Yiq+WjzmK166PUxV3RpxaWG5YRe+KWRjfRgVUFkxKfV3f6Pe
zNp32D8LNLfhz21OsJkmfSHLG+AWQbZQ9ERg2Jfp/c/N9YI9vkSgRJSkipYnmk6R5OgnSOqaKFq5
P/e+1ibBzS8Kuf6AzabEgA/3JESqxRV1KhlieTuzzJC2gJ2riejDOwDTXbuvpWHYuWHQrsACqC5r
mjmBFDSBaCio9HJpQb8+Vltfi5B1lb4V6SB877irgC6lsPDGhyJi0ByVmWKancFSZ5VpyhsGIh8x
38LH+L5mL6AteoN40O5/9BsI0hDE/KZiQTExYeZdISkHqdrn5/dU7odCDds34njbxS75/zyMPCen
rPVlRE/BBiVYpXRVoa6OowsWgaKZeD/sRXsa5srlqhDIW5Ox7G23hkJzLHy4zAPcstVZc5s0QMLb
XYwQVYidXv7+0VrZ03Poh6XN8/DF0prVhYsVcD4RMIQAh5sAtgG/8lT5axPJ8mXumSZv+f84YmU/
Qnd5h+eGk4XKvsvL5eQKFTnywW0quZbUsq0lDn6DfCsu2WBM745n8xOnUoWlpYs9p7cZESyOpbLR
tE9QlBOlbWqN+5wGChAlxx0tf6KJAD+fvKt5JdsfPPdMgH9tMVk/pteAcwa1zbE87/oFobFOuGni
xqeG4rhKh6YCg+gBRwjizD/Dmn3x4EA8eZtuWkUqNrplmxBP25990Dp2e4MZP38MwRSORrYrD0hu
JjPziwxZOtgdg9wzcTliB78zmDdf/iqAYn5vDAgg3XqT9prLlq9nmxI6FbdFK0OSWH28Un2MYWvn
Hm5WLQ4UAP44jv3+WmxtIVVmcFEVe1v8YSS+65YW+mKTiL/QG8mw7uLYQLKu6OJPa+gx0ugK4dIR
tNq5QJb8sk91AOvuFOlOrtNWg9WbCOtVUmrfUTJKkHFoRaph43ZZGCpqQdaWv3TTAH3cvv/8mfB0
WJU2QeyTrmlhNLkGgyF50VR9GPpftBCNyYHdeAiMmKU6hXDYBKG8YOtPA7BGDc7rp02VinGq/fmG
MnvoEF5+jAwsFbJwCNd7ckfBHhYXZXJggO81nSQ4ajfAWWfdN27Rx1vvhE9SNQ9VJaK9EBZuOTte
QjSxr71Pz3y+NpEnq9ZNsxQU40RBzMGjj9+AkMyy0n4lLwNXI2h+l4YIlFop9NqbmymprfIhQCvV
GlxRRc1iqh7zsDVoIrVe/m1z32O1m950Yj6TcmXnAxDkuYxCNYU9a3W0ZhMFwsA3nhSL+zHdX9lN
3fQC8sKPl3Mo+yWfba7oNh7Dgb4fdVhbKNlJ1yaawSoslZB+VTryqu5ChgZQAiRF37VgiAc6zQze
lF2l6px/TQEYH3Fodjfk69YjDNUy0Af+WPxYe3xqhQ7TJ9JInDfY3CTtksKi8WsINX0nHdrw4rLr
Q5nJUBhki74u9UVioaM7g50Epa9qmdjb7mZfU90J+tMEXQMEgOhZ1LST7YeZme4OU8Z6oZgaimp2
el7sugtHQbVximdY0Q94fsE5nF5R0U9E788vjHhi/LBV/hFqP9UNyFgqMnCLGVf+T2m/axT4sNbW
juh0JZHBBzh8FGunvzamKxUR/twYk9z97LWX6p3JXWz2vlfI6zsXE/90QsnZsRYpHNiRKQQ/4F0D
sG4jnxsH7O3dPugHcXuds3L//MzkCZbFq2h/RJirrUHyhlz+cTQX2Ze0T49x9GfIDIKsfPZPt7Zs
wcuR7xh0x48Qaw0TZGF9t9eV0dEBHSUjpv1Qqt954J1V57yWe9I+ZIYN9slCNy3ZuRMCtc4y0419
ABToPXdGETPdBuM1Kwe9JvuZgJJs+GKGPvc37abH3L97lg52c01sItHkeoOGe3ImQ4xGkWQrDfmh
UJIAHSsZNmhRu43gTJ8gXx9QRUWeB+SHWuYbSaGZ2awNTeR4JCRtPghm+xPZEidPVSJ3E/mftYCS
HXFUgLNEImaOHaIuu7o1Pu8FjnUVEKtuH8f70tJz4Lmv95wiXDxlWadTZ12usmjRK3aMR7kCzlrz
rQ8uw1sYpRHIF+po/rgxf5lnpmsUnSC3cMOZ6T/aOAuoVD8/+8MHCLc5M7afnnCLLZ7F5vddx6pP
5CfyidetRrneBE2yodL+ZvyZZrCWr1UTPAWLcbvX3P5StYei8RgjDuiWaCXWLXL9AaPKIUaXXz2b
GFmXTsaVwNVv57chj3TZvBw+BkKDbiuJaGoUYG4WieztjPzrYO3N2N9x8VQ1FaLIjltRfWHhZ/R7
uVnVWvca9Ohk4GKL2FPxU533UnrAQ3hRs32IgbrWjuqHQ2UogO6TTCzczf3B++GpRBAT/BK1n79i
xXjTNpPd21OQ4tco881hMsTouCYHJWWonCk9s4qhFqvONK5uMFgcJbXTGdzsn24aZQtwFqWs8m+J
C2W1n+VA74bXLHX2aXGBia8tipmO+P+cUi+de7A+5ufNerNqUfTcOXbP4+XhgsYJM5Hf9yxUAwnY
pxdBvHaTm9B/Fie+9s/VkpbWAimGo0Sq+027GDHck32o8tts4A/VkmGh1acD51QdbI2HX2TWgZVF
U/U8zVRmloZrSPzl3E3bRcNjofYAMHoJqBjs55VtuMwnBFp2EI4M9veDgXTXrR55bIoFpVQMwxSn
cUh2x7garh+xDgg2wndhXobf3fd0uWpnF04IBs26XocWrUXTjWkd8vuqh3dzlJVLoKPMyt0l0eXA
vGs5Y/5iNMNsC4HyKyIaQQGzxAgiUPWmTqhMOom5Dh/jtGu6we9+uJs6IMnPPwJKWjVCRwyzkiM/
Zp4aq8D47W0dTzask6sLHkKVWtTTHJcbTkpkl5MMZIFsbY44KbucCC+XrGt71EqnRU6Vjrbuss+U
wYfez9eyi5JMfgl1ou2qMaKTDZQeR3jS2mXrRU5bvWm/sASadxjCEeEXT4YzcR58/yvXM6Qcwd4L
6tp8sSYzbrWbV0UNQXaJqmPYtw5VEBilJr5qa/uAYmZjy2oUi4SM3uxlzob0NpHW4F/1cQSWbub1
lLxHQqbPDRF7OIF0dUthudDc3YaUy/MH+hT2vObSjJ5mKpljg7ZRvFTMtmNrKSa4O9CRA/Fo4Vuo
go1H3r910V1rl0czLOapV0ijOtqAQN4DrI9oM1UVEC4KghighwNoTaeIr8EAdANi3crJtWN2mHCO
3TpYf3FBYMGDE0Q98POq/UPK8NxJI4jT3pHkfJF5UzXS8Yp9gt+b3JZQDTXNIw5ejLCo03K8XSVZ
396+FsEkVi7YgqTLOWE6eSEWPxiH2sDmFtHT6tW3jRkPWWQ841zJIRVd54yZnqOJ8qC1dLR+ATDt
3USep/Y1epw0McbyQ8XeH+G3UdT/zHg2as04/JebGLz9auzPev7hTbqQRXOvBqpnmVFdZv7yY+AG
UDk5GPhzPbCq1ElCn5NeYbsXDoF72CMMlWaGOjMPxK0Lu7BQL5GJFov8tqzHbl6pWw7i1Ib9Gkdd
EAsISnpnDOAgarCU6Fq541myq9szYirk1mrTiowv3ceUK++ILqo7ZNXeG8uMNZF143xtNmcoN4xy
bmRRG/7sVJnZVbQMAYJzPRmIjaa8r8bhRIsWiNWvbokp1YysjGAvQi/soDhnANzS7iVmZy+3rhUt
RPWlCLYmqjc7l31abFOsel144qc9FAt8WDK1n0hTRFiRlJPU1sWb1eZXhOel/CaS++AluAxJwYIz
Snhhchy09DIzqyVUNo7njG/aMpIRhETwIORPXhd+XxICzU5a68da3A9V3ssOrrH2pYoiOL2bndQQ
bRwFxczZjYAxTWyepeQLyH6BM4rp6HsgXk/Lqq3/R58JsPC5CUd97EgSgitdAUMYTmu0/XpWCbkJ
b/1Hy2U2/tDlz2mI92ru6QBNG4y6KKCvd87I2XQRMU1G4TweXcsmR4TPfsCtlpiBqwA6H/FVkKbn
Kq/pdhNaLoWMnkEydXSapami10ZA7/wiMt+DBbFaXRPxh9A69zpjQs3pL+wj9GqWVX/onB2H1tol
/qHbirDnTc1ZGDpXX0mqn4+9XAZIKH+dWZ79Ni3CoKbXEpmrrRm+7GApSfR0UNIHvdqywJ951CQY
hn966fNaetdOTZLy/rr1lFQTL8FAuVFTYYYNmqATiymlpEcrtGTfsxdmUi73cBwLeQSInsd6SsIQ
PrmuTixtftuRB5RanQ+UA0ohDKeqZR7ml7rpF8w9BIqaYzbkaDXRuploNwWRxaKhbN3AtPx34veJ
bALd8ECIKNlKTUXIXmCtv5SCPKvlnB9dd1JEyDd/xJbBQ/RtoiL6hjmVgWf1sLXT9avbRfGK114Q
Wyz/RxYdLZJ96YUs4Z3ARGjp70IKB6gAfwJdmjoVegoLQZ609X/Lw/2bQu4umf5cCNsMzgd3iI9j
Y2K6T37UHOr/t04xNNfZTwCjHCpyjT6FC3ekH73REGzRMjqt+bIRTN+y//bsiKOebuByW8CV4C2Q
GfIgJjosODsqsqgV0Si1+eCG48MjqPpTncODJf9YcpU846brf7Kfbzo+Kuv6UolRIy6VAAbpOttF
r+9lvATJXFenapV57wREvXMPi3I0zrl9EiuNqeiVXeSWVf76MqtFOpDKMNo2CHM+MvoMlR0Xnl3z
DR17Kd2WWDCChhclL6ejoSxC2jEmGt1IembyensmSHaEqeswrtm9+5I9alTcfd/KyjVmoLXPnBDB
DXwOUvz6GDw2y/T/UiOFHpM6yf9bXIrkDuqpXDM68tIHJsBtqonEwpu53K8ochK7R7Jg6rNmLo9F
yKInIPS8hG6EPiTvA0r18M74URy0urY26mozkK4R1z9w6HEp9WaSPiILjiUNV3Fi914MT0JTJAqC
9qPnVWTChD+amOTt52/2eVw2JhoaNaJ2QwqFEJxLbV08k0alPhqmdCWgIQZHOOvM9rwuGN1UJG5a
R1xH7KTMhdjleClsNCl0kHwkU3MSQ2x/RBluaG9ehs+RCn1d1u52CKKZuAcvlh0K7mT3yS+auUtv
zMZihso+ZQ/WADmeBq//Rg8M1SQYHGtevYZn+LRin2owgvJNL9i76o256zEv7sUbY0zVF5xWJvCj
n4V32AaAATqnC475e9Pm/b0qvCMgxHBC8rXq8fBT7L4ynxGNXfIdNPCNqP8DOXegrGQqk6YECJsn
AS0QnnpEQi3+7l9n9GbooHoJzii4xtGo+HaZtXZuUVZRrDiBpFOHgVyRlyUVvIiEO2jZN65ma4B8
vGQR0RnHPL5lgCYTRJOY/JP+1aVW3lID/P2S5+5fhHiq/blxkioAvFoHwHnFgrMJghEpsEphkPBk
XDNUA6/dGGg4RBz59YbK3NxgeqFNYQYpunBXlafeFp70v1Hy9/VhtBGphg8DWCdfp2MH7vx/1lTv
XdHS2ViZDvyAmbTsSlQc4zQndxbaK+IA51CPCquGLqW7VmXsQqD32Hwn2OnAWkXbMClcLD2b/EKq
ZTezN5GQvwL2qaanjid6cCBVeqU3l2DlE9wTSwFE0hsyeBBcK8e0AFprv6+Fraeh1UgHGdhVldm5
Mnczwj5DxsfLQgvLJwT2cQT5YhOMENEwUkGMJh97QTREpCmox1evmLrWRbLUGGJvZCRNy2hJKyNi
2nJf53CsvXwMnLUpjXAGx1tMTl/QIDbsEFrxYZf2Ksa9to6zu8wz0iwAAFUeG4ut5eYAHrk2IPUp
NfCR+YgHZgEryYi8M8xFxHvTg9AVMtApf4IXw51RvU8h9n6zfPtBUVQW7a/+oZ9R42m6Xz/3j0D4
4gyKMvTo+AlwEvIYYz/rhpQLPA8X+u0nibukCE5WlaVl+Hf09gHW8mydv5TqfflwOC1sPB9ogmGv
MIgoAcEWA/zi5DgsX66RGa8/Kh37JKqvsdj7PYUrdUWxvB7oY9Fc9Rv4oyUvXcJHuSd69pqaxB0b
g1tyYZ4S4Zf3c5KBg8DVRZWYeKm1Mvr2jXvXi99HJVxt1PUcbzWSVKJMVD+DqnuewybM/e6IPyXO
+vH9vy9VCJWLC8u+g37kb4U4QfA7+kZAIGJpN5WNOjhZUkqBfYvHiBu/eFpp8e2l4lwK0Th0420O
mQuw/vPPM7JVdJpETKarWSjneLknu2ahMNgpZiVh3uTy+2mdg0YucMFOzt1zxl4QMi8zZcCd6Xti
isJsdJTGXnMreOX/TWIWFSFZr0ZY8OSdPUSYWXgVEOJ5iXftN2vG2gEqwwiOiAUGsZ2T48SiCFzR
dSPsJ2QC3i4HmtTD5g3M7scq2GRWMS1WWG8d//wdT0Vuji3w10j+1oEUMJ5xK4io2mQAFQYICff0
qZ3ST55ASn6HLYFmTVZcpfszgM369IDN0GK051si5tIT2Mdjhc6GfAz/qQcC9WKZRV4FNJPuwDzK
RHTPsmG15RkUZaXuNct2qYgatG9c1HTp8cyNhO59c1oHKMDaaGPjnxVFqPqMfXnh0U5+ec+DMNhS
aUQxDUxOP0yJbXtjjjipjMh9fQIoqRcxum1XzEFohJcYgNmF7rz7xIWodtQCwt806BzyYKGfqsa8
LLMUG3v3YP3nNsq6Mlg0QzBSaIBB2y2vJEiHrdGPXp/Y/JP3jm2Z7fLoVJqBY3hxs9tL/aY9DDn1
DrH1yQUtYlei6nzoGNwDgTxeM4OyQtAO1bqUTK2dYbkB6tRVOyzW7N14VEifiVnH9NBeKTeW0xZY
VbnkBleVOYClCKfPNH+A1SlGPipe4kDbVoOMWettuUsi/mUnKwnZME2sLEiXAvuntDSIY3MLzktu
Z8e9IQroI6qc4axNkOqdOYOec9Np9jUrouwp9aCY1RZLsmK63V9oHUs8Opu9gLwsrni5F5jv6TAQ
zbguGesIeYwnsFAmHuY8UPvQhJ/DtZ/Z45+cqxkMJzXW5YITtR0rwxi9p4tCRMRNb32Ndxb1BMIP
8kuS2o4ZQuNG5ZiI8GwEyYd9Wc+647vpMluokARaiRhI4mYS5il6JYKkHzgpApRcVunVfj8LqwtM
UhrSABT9xA1PlUj/2CzsSpvUeouxbsHGyE1ISUeciD+6GaUQYxvIjU8sxMpFAR2wfK+G60ASTz44
+TOqJhPH4ZpEb9y2cr1qMxzcbgZmu9bXE7hFRfJ9c2yanNEy4gY7HZto3XQGFrFdIZDSiw4G65Cb
4fQEsO6I9OHX8LEZsqEzfGJEcdIm9koChdOX2O08/jDrmBJjwisoVkzecIBCIl9cX7PuVgVebQvR
s3flYzDlpyoM4XJfXxeFECMfWrzYrW9qH5b+tua9jT3M12PXKpcx2RHbl+OBf1TBdkkM+YuWnHXs
4qTa67/NheFE3s7MOK+vv+egphz/2uSI0Cmg2GhnscqQwSrczIL6CBMh2b5oI4saC94p32lzV21L
07xRIW7+iRUDRPXvwwryYCi1VpYCfbnY8iyf3T3zvAGH9EtLABPYxLGcQiUVfEyKexPrZJt/o8qr
cCl0CoA33+dpxapcPRKqGSVrNDMCgS0W+0thZx6L8kFvfRot8typ9qP3G3l19ciRBEWMz1zU3oFv
TZDaal+HRe3tjRPdFwYCWftn75i66BXgj2w6rSquxrVAsBcGtKpWXWmnBKlvXMYo3lZOwvzAAKm6
cjRYSOi5NaBFds+TWaQBoQPRZ3N2aPRoXcnmBBzdBnTBVDLwGj0DTNEKrfUxQ0dZNx7y+e2vvng+
1YN1ksIxmI4hpfy4dHEkfujOn2d6uvdJWz6g9WYg/sjJvNZXwyzU9HnTKI1rjEj46J8arFHzy7NO
dlf9sYr/ma40Kr0cplACe8BUDRdO5Ne0TiA9fvDkSXoVB8MbopyB2opCpJTMoD3oQBTYx8t/1DEp
Gh0MFlppmBIpjpYIhxekrNXAdndOin38VgCVYu5cYOOw2zFR/4wS90wlSHBgiQmloc5ZWGz+Nye/
KxfJSyMjj2hZ6DaoWYYvoQ5VD4gudQNGKk/bQdce/q609Eerc/qBkE5pY+ZoTtTORafImZrQuPxw
lPPWsDoOwaXVDD5xdIzVg4UF4KoZzkKQ8a0x1PUuxWxgnbcKtri0ht0NAahVwppCvCU2mpn0WcoT
OCrjGE6yspR/NChggjxPLxS3r/tjUXkOjmXGjw/b8A6GmLSlw1HXpe1nRnbLAPs0q4KeATkYw+0L
p3NMZcxezsTrgYVIuDWogrn1atKuKCtZxWIu1Fehn0k/VzrYU07eJqkrap0ofRl+3pHyHzjXDH3b
kneljdo5IRh8WjL09dauh3HdlEhlnqmYQ6o5qVL4Tn/kk6Ze+mzCBxNrOHkciDJLaVkNwX3bevqp
k3Cdo96bq/B3fU71XSSGLZceZOt9gyBBkoDm7IbmrNpdJOz3a/otbKPm3NXFMSTXmUEV77zQuC6+
va4Rj/e/PqWQFZfLsa1dzv7m0lzx12KZ3ImhKE9Qz5zseUPon2yarFn1tx3THppX3QxO7hYVot1B
VmfM/+Jo9yam46e0dsS6mUV74TJLHaRenVkcCMPjt+rBtPIPQ3D8Bghpm0QiFiJth8hmDAPJj8ks
lu9n7QpwW8bfQaDXGHMSLfuUI+zy0zw/qaunnOBNXDY2HhFqJKEM1Dmf+KIQQmeeQ1ia0c+UAkkD
AGSzTMEwa6tCtYe4gIF8AoX+npQTpuzkR9MZJkBsNFjyTBjeoiZFA0KV8XWuD5hQSzor/8Wx287E
/I4b0bcYtCydSmVBl0HSw+YUbfSKLRvHQb5iRKTFR7JnbSlhS78f8UlrDOP+Fv6zYecPJWCM6gYv
NV/xwBb09HE7kEZg0plC7xGoxn99AlewESCMeirOPDxz+4a8tToK+IlRdDoqdInQeUKi0giHxnEH
v1n4xFik7ayTTrJ7ijrdWO8w7rKcwel8MgTcRhFH8026gavulwt8WmkM2YJRhkQR8VPQBLGTvmc3
GqJKtF2xt+T5tWajFFhj6c+UgHiNajoYbuLMy2vigwEXhw8lO9eFd933rayC6yZ2PR0mJwvyAwqZ
MVNut0JKl0Nk02DBEyqW3KhDG+roAqQFfOpGChl1LkJw89/7j6zKF505b+6hiXl0GE+u96i5jmtn
wk0KDMSQGsgX28qq9r6zNgOTOmcX1jIDMRkfmE4o1iQNVY1BO+H7l1nC12Z/6mXw12sBXC/xArcs
RgwKsLpYM3WYMf/n70g0k165EHi1Iy1t5QrZRGYiEMUlH9iBqJn69tKwzYu+0Gvuwdx1E31E4vRj
rKGNNd3Tf0rGNpLOr3is0xef330X7U6z88vqgfYxdTvxSIekXpHeqtmjE8fBG3o9t2uVna2v1Mwo
LeorO0SLab2p54YCmtTAptI/pApgDSTZC5xYtfGpDgVOruNkgNrC3iwj2kuTx4anKD0xUMnHvMXu
690nolag7xYS/0mjLa+W3iX+dJl3OP1Q50exHMp5PO4QrA/dYFtnyeTmKWd4noY2QNvhP7bgcJDB
PQq92gbrvAkJb6jhvyhthFewUk4QoXsDl7wVy9BKw4PBZOwxm3Qq1o/7HrgM//iVX0NdjYahiJAV
3WBSurdCg423lERftDfrVrLws+QDADNV5wxtE7Q4K/IIQYBf8193f+a4jVTlkOnY7sLvTb/vnnM+
fCzrL4cM6rK83Msui//OKEEsEWaiEe1ONzOBtpdkJcJZExI0fd6ht7xg9vjXfZSWIQuGKaMuaWJc
scVQ4OENK5oUvdDCxZWGoYdAQ6UEqWOHEp1Tefw9dLa/peigRtorRKRnn/N0903vxv3NDRp5bDRp
OQNpdTfUe1iDhkcOEb1d8EUWn7wSj9wCLGJ81Fbw5xLccSt1nbG/KR2lQh83E5EU8UwhiaBFGbh8
9kAIGHtal0rsJ/nBXh6XD8kaNHk+F/3IIPsfu68XKf/HxqRRRsP94UqZScKH+wOq76miOJQOSl1/
1QO0v4dPoyRkds5Q0rjK/yNLSdIa1uUv/nmdgfKjP5pXUYtjh1YAT5xzHb/NMuBlKuCnVHIpyvnk
3gQ7iXWnENaRtX63Cb1NmTAr3XSf1AF1TyOGa3y1huQrKhSpVmse8MApme8A/rHd2b+NIX9XYG1R
IWpweca7nhuvrco6L+WIpvDertXwIq4QRd2EnzbnHL8nIBw5PdF9LWbE3DYiAKM4CUkchyFbWURr
yyoW20+u3iIeN8B0midYATF7D3bCBIMQ8BWfnnOxmFvV9La4fG5yysNtucchM7ozhUoN9EbH8dgG
MP1Wv4mxioQzkVeeAJukWmluWL4J65M27o8DQ4Bq9C51nfcqVTbK77nqIvM2Uj0K7m6jxlVzXBUA
0Bb56IfyQkSeiMwuCNccM2si0TA15zEDAAt+aQH6pid5s3VXQv+88r/54s1JndZHCELzhxokL09W
x2FV8bV1VAlwe3zizc2VZZIbxsqGQBKCgw1rOOHWgvU2QCvmh64Ljj7u6yBKF6ccXCdIXwTCLocR
SAZQ4eXp5le5UpvtZi4Ykgr/3wpfsCW4A2ueI3K/kXTTs/R2bNXbUvz+ptPtT9D09bBerCIuLzAI
pA5Nro3Cj4fNXIoOR/K82N7nv0wPJ4RBL7nqa7gedCcNIRSwP4s+kx8DCYXcmNJkhEXi4BHEbHyz
ZLxCppdgq3mNRyyJlpn/y3SUCYn4VqW2MDXvtCfUQHGI3C69MbXS0O7u1+zirkU8dGq5e2XstEPD
/RAru2YgTM/YJHgSOD+MGfHw1K1EXIvlLCoAsiPKWPTHUuf5YUOvw9nP0GCsCaCxUaDcDbkJLdRM
P4qsbaaNwBqE2Z/nyv1y0Ka90/vd/aE1RQr2v4kzNNneOD5lcKRsey02cz78zA7vBpghP9iMog44
oFh0m1SwOkUGQ61lHVYDW9EUhifx4fj7v8bd2RXrMk2HBnJv/na5NQn2rk025LJuzepVKOs/Ku0m
VxkV+Sz2oU4769x+/6f3rZIp251pohLkyT1unsTA77bqUCdzm9Jy9layJPhJoOmSnx/hA+SIuXhN
uDttFhsIf692bafewZU4zujtnSfNJtQl/WlPQkquyeU1mqD0pJLG031VK9YUk96Kbf5Ir2xIQAGt
2bHRqJ1q8c5WS8etMeQD4uL2jRFxxB1a/PdbL9TM4cgtt8m5L4zKnsU8oQGxJ2+hzOp0hHqtZBSo
ECWa/FSMrLVOwBzGGVLGcZhPlPW4lhx9pxH9PwWUHkC8YWn/M/chgRjyW6BwHebFaB7HmxY2FlZp
QXrHElz3Br1uVOunkkfF+wk0r/cQrwExIRvbzZdvtDUv3Rk1N+PV6ZA8PQ260apCcMzhGaBnuISl
4oI+1bLmpAlP2hYhQcfwa8cngfPE0kmA1+Q8bKgTsVt0NLLlb1oCxL5if2bq4CVVv+9ZPHRwocdV
poFFjukw/ZQC6pMnE/y4nJM6REyhAfu4DgoFzR0rwu34+3MTUmPIf0ZBpqx3pITqHomRfp6DyuH7
OX9zmxIBmGV5DyYFX9sz987iRD7z2evyrvmIuo4AF0YkGRd0l5X4o3u8QfZKrVcEtIAH6uocXSJt
RYvrl+6oMw/LdPbifa0/rSlAWnhpERV58fYPEUnCf0z76KWrRc7uYghvet+wa1yjJFuz2hWAd6dF
mXRm2DDJ8oUNx6ZCiAhUyNryoM7u+t557ICb3sOR4Ab61NNg5hh2VCvkOXP8x3Cm9aXwQXVbUF1b
sdyXfTye59WTIx/4SEBEjbDVX/Pf0DdZ21nLpYAYL49QmfgBz+dBIaoVl1OnHjeOnh/VUHJV3/Y/
Ss25sno1gi6ztT2bOILZS+l2nSSi1NL0R5PB/v8p11EItfsO4uW+ZbYuKpsGLjgQ2Sn7RyBlMnmZ
SMqB3PsGISifo5DlWH9yGRZ9Z3VdynJjWUH0LPhCgNM3Cs7QRDSo3+ISioRfScZFvsXxyNgwyIVV
5SA8UPuCNV5TqdsowCC3OrQe/fES15u69nANhXaSdwkFHlgkCQ/eu55eyE/lRaxu9v3E78JpJBtW
eo4QJcnn4j4MHg9e9a0R17rar10U0JZ7q2AB6EFIZFTlQaL1kDUCL6x/GOUiguhSOSE6sTyMWBOm
WQMS+pC/mW2E33v8Gv1SlHMvZqXygyMvI9pc+kWxdOJlLzgQdIKcbFIDzSA6/Erva+IuI0cf1beP
DUl+wwSWo0SnbVBV1MESn/0U4eGKfIi9VS731ox5LK0n8soimxM825KGRLVd5/qADjYC3en2NTtf
KhCQ9ZJVdB/4gl4nuXDikiphyEt4GaVeTMbXShVBMOPsj7/nymmFkQzQw84sCGrUJ1pBXh6J5tvs
2ePEiQubYOTMiUUcsW2hXQQlG5iMw+QQDSeQQCgXqCdcHY8CQKBAeyD0Y6n2EWI+qjsf4eoQi+P+
rzAcsV48C5eI3eCURPYlmHV8h1sgBynV+Cbx/CoG0p4CagIdtTiNo4Y7ulQLiI5XoYpp03a1QLWJ
0oV4yprdVKtKB2CUQSMaqN4fAbo5FwxHaEy8CsRd2ShKq9Dril5XXJPUkKo9PKrC8JP8TAqZHlhm
PcUv86Fnw8lyCt93mXAKXzhLaUkFXxxkfzCBLbukPoPdsmcqSPYfzg/2agW2uL8QZQylVuIY2WEM
VKLUfAWy1OrsfrP3UG43dkX85Bs9jinY/V1I3Aag3aAmLp9PANec2ZbLiI0rR64CAjkvRvITVLrA
SCZVZOXFO1etLDzux0j/Qt6nOUnkuI5eQxYQv0SIb+SBXHzKFqQ4YEidZfQrsA/jeDywlIo3WAid
CJyA+FqNik5q1qKB8Nn/dcsQQPGf9vnY0kfaHeLKKUdSvwwwUuCS8lVIAQDN4LbhL1euopjUVV0p
vYtp2K7zd0YZNcBEjBzDav+9JFlDi9+6s5ZS3g6nDrs6B1hIbt4Dfqlicq7JgJOrWZm2UScwap2A
hQJqMyelPknXp9EDvzRQ8XhWj6B8OhsD2HvzE2UFUuEvZqz25HbKIoY97TVsO//ysF+4xhT1FfVC
3MfgErp4+V8w64hUo5sya8scjWSXxFabPJA/g/+gAkbgniTFnSrYykPZi13qt5BplZSmsm1XeA8r
lUvgk5PfbmO8Zez84Qo4ULkv8GzvL5yrIeoD8sh8rnhZGczft+cbr4vauBIEhUQzj4Iggq5zGDnz
v8PoJ6T5mGxHirLLicw4lPCl6UjPsfR1hZ+bEmwO1HjL4lgDeHUgV2DiGQUOIYKTef210aWaitEj
WZ3cEzZ1rK1sOm4XPZm1HYKQgGg88dT2YsfsrV4RDw4QF/KLTqKR2t0vtqk/x8LTMOYS4lHNdcDq
M8R7wHDXiOcNY4U7s2vpDG9suvzJiruHhEVNEtplRrUOAmetxdtOS6f5jkEz5Q+tBqDuHBFx0QF0
w2vyHppwVmLAXzBysIQuyugMU+opYXA1Z4Jjuj09WqWC2TmGSQVDUtkpJyGrvmfIGh4c2O3bIhr1
EER/e4tAGYG2mLrNaqheetQsaxdzuH1n+P9ZFXdr2N+lVmmPFyZYCDPrV5R6/6R7LfWOc/w6EPiH
URgI8sVRc7sAp/DRWQ2o8+7NK7BDlfZS6f8BOrb44Qn7EmBl37/8LHP2A1xWAOITk4Eb5iB4AjwW
io+OSFyCcjq7/+sfGTJ4XdbSBXaBdHt4JCzFXEqbF481GDHE2mhNd6hHT1gynrr8KDaS1WjBKtUf
v7G6Ba7jOUASwDHNdJaDOS51psMr7npnvpWCscAgvyM9Dn2bbIMovuOwCezSdNQC/+BgnXJHQt4A
q39aUYnXlOEvS1qpSrEFxUU3FgGDnXCn4ckwLWYMzS3z5T0kYxrG9VQ2gujJjriiY70lavievCT+
rA+AFjLIy6Zj1lsbnAnzLw4UDkatrE4e3Go7JjVpQOojKGfsCrx3Slq03qP1kqWSdzxTgkGQdX08
q71NVSEiE/1YoJK8aKxn2DMhx3tQUkXHxEtsXdhWuy/l6pYOpkj/GGrRpBlQnIXX6peu0uSmhX6u
Ssedex5TUNb4gyKq+DzQnKIVD7yw/9MHq3CL8Nq4bg42h2/Z7HHuM2X/zwE9aM1ZxL8/epqcD5Fn
etnSJ4lSVFo4Sp3t8b6zzoo7ZLm+0lBBMfXZbRFjsxWFhN81RRAtOMGAY0GKbv9zFpfjY4tVYlt+
K00zxp/8RCq+g/rpljqshKMGNWLLlSeu4mhF+CX/XeJHT+g4zyAXeKMJUHLYIB3quMbPpMNs1yu2
0NrDuyO2uAPyqWXw8PCmQUYrbF/67BHBak5OiwSwFooowsImyU0zTU8BxIymQNSTufgPaDQBbr9T
Dm8LKuvAZLn1UnAS66q7WrjN3oIUaklVEmjq8YgXZ+/zwWiIg/l+ou9Z1Qg7MvJ6OkL/f+sTWtpt
pqiU575hQIkkn2fwli2H2iwX/3Ra2zljmjkceiRPZfPn6eHKISxrP08G2+kQf3iX3syV+oYg4WIt
KVgpspOBWlEWayKEoy5EKtwqqrp6bMlqp1UERIn8Wlydjdtbul20vwhLcbP+Ebmp04UZXWTxORnk
7af4xCMCChER/BnRagAd7Lzc8C0xkmUHvug7+Xt0WxAmqe7kkdg55Dm6b7in4Ogc2T00/3SkxYHP
trysZ8aBubhSLXpfFQ1RFEcrNt5IafHAWCUlceipacF4F4CFCPKDBH5OutqzH7mKQayakDol9YTA
GH0Cd3Y3zLCqE7NU6kK4hLtvQSw5elQibnNvNXr+SMir3UlTXtb1NFdqH5bqzSZegrUfq5zids1s
XNfci6x7SIYGAt2yfWIMYL7NX5ibj1U+bUH+jXqZ85G165UGbdZWwscX+ksWXQxSIgzK1Md0wZpE
YEojqfEDYxB8w6q1gQiN3JbkNfuT5fIVkchZZGIHgb5DSN/UKJXqxP2MKZ+YBnRTMNRF9q/O9/C7
j4w8+F6psg8lTMoIxOwTtjmSEvdjnu7tkjEAmpKwsVStBEUksSSKGpP/p1XnYK3SAwq8M4L7Teeu
yU0/O05rgcKpomtxjOQy4gOczPkzTxOWnEZCG6ZpDucDKFPrh+o5A5rscUxvnwZMp/GOo2vRxES3
6zzqcedFNOF9x9nrNmx090g9IhfR6E0GejZmW7jVseFAQWCGA7LtLfsXIpHJLgg5mkzDIFcOethY
6xGPIBWDck4l40EDDnBhia/MoB2GNUvYWHhsUwT5Y3TkFD+CPY+Yo6FbRevJQYHvWq5kBt+lJ6W8
cftaiH1/g9Is7TQsv6YLTx+cJPZrvgt31GabiYU7frXhRhLKG8A1CaZb+s054MH1Ps6C6S0HLfl4
d97++IoLEY3cNSQy4CDHdJ7lho4Y6zhNlG8bsJq+/8615nHvpIwi8g25uBZCym20vh7/dK4Z37MT
ESEOxnzeUEB0lG48IJL4c49gQkbgVq9o7Jx+ddAsICU2JyLePTnvz+Btrzce1wEPDCXIxg7Zws/4
Uu6lxJPetE64wpl7ow6QxHFJ65EaljivpG/QCiGCVpkPT9AUsxG1Hc1nVjlSEJJ9cWlAhSBVZ/qs
Lj/uCj8juhE7ohZ5Dd9ZkZTREph1XSah2GxLlt8JjG+u6va3a3E3JAqJQPMxJNR538h0O7gKxPu9
Otr/axdJi3XODqUgIdAvcPb8hyATNDsR3cQ9jT/t4jy32H8CY46v7DhbNFKRdh63VcPVE+EHVCt5
vZzSMUWJ3eWW7n+Dr1hJ61QmhVDsX/WDYKpgjr2WdZzmENTMsSHdBNNZtOrW7uAaETiYopi3xLmR
3TA1IYrZtgnPx5unvsz4aA3M8bPpSNL0KuwgRqi0aBNajrFcxZKg5mK/IfgEX1Znz7/2y27mK68k
Jso+wum7aHtWA9S/nLLBido3QFtKFGrljZvnxet/QExyeJ3kYRIvP6s0nEwqy3AknSA1+hM7SKQH
G1imd8sGzQ25xRHa+r2+/MsMteEWZ6A8bieG2GR5J9MFl78xB4Bqe/CfZg4i8LZ5ylN/WkuMZhec
BIoB2jC6Wnc1390Fy4pcCHN3ob7RqnXWHsZPSpbqtTfaxq6GvqgMpBvkJg8rOCi7wDHDJ1wwJatF
k9TyqLBvOLu+Ni6ARM3H1EENNP8c94D+SD4GG8AOOSNw8sUB2k2M/707MMXoXUR7S7aScoVSrhXx
V+56z/sujGHfYBaVXVWDdwmU0zP9A/gOfHp1TFaSTntFvWWgKvHtYC0q2NWcpMi+Y/HPWxWJ4irw
7vOa1Ddrai0xtMRGUJh40WGY/ktRnOML9iWQXbYZsyNRqefMrinImvQnpuvwrtnmS8V9LMHMh6LX
jO0lMI6Wfx0A1kmHB3pz+f4vsJnsxXwkPRzkmFT0u4r47H4PoxswZ/S94sGYZT5M7sN/JGHeR2Ro
vIAaj1XDhA/UoG4RN4Yvu8xKP5YpIWJlAZmM2qiyXXZ1fafLJRCyb+v9F1gXq27TUj1uLWxjU8e6
PWuv0TRr5og9ePeKQSJpKCp311h7NAyG28GR1uJ6p10DkXzV4WafpzrG86ZxN3GNCrEH6L548n0k
aK1NlVxu2qe2D3dQjEQLbUl3r+kb5UctzJTLLKQnjm0wRK8W0xehdm75YIdzim38dXTA7CvPeIRB
pQD12bBSXW/SEcbF+cGcYMbXT3otMwQkqScaCeLMQQDwV7tmyZj61H6D/XkV5I7kEdOU9QLu4Beg
w0xNGCjlMnal5qPFuhG0ziTmjtVOoxgO2Xw7oyDca4p+NM8QlD9rPmmbUdQdwAUmpxoVCX17fEI0
ESgbNOYC2Eb37TxQHSoUMZvKcJV8iWLWRCdoMr+T/+GsrmkyTP9lhyd5SJdZauSlc5BJ1RR51Ory
Ya9KQ+dQ8b8UAonloh836AUwymNNfUqUve0nEbtOH1YyK8B6BMoI3CDUgRFTnZSFzOfw0FA+qegA
LhOLqpyvcvwaW74KBn6/jPOuoU9Jgx5K/DCwLjPnSyA2FGAngRD356Cs2Sp/tBc/rowAxobRsAch
oNrRS9ePRxmoU7Q+56i+S8ond44GE8nCvd0RJ0+7HEKvIfzWc1LSXoaSonNrJT0BtuKsZG1pQKPJ
Ra4+zKeuDOpCOLkkBpdNu7ptsLU7ejOePaaDj9CDCi25Xv59ORpn9u/eaVuCC1zwLIyMgeSX/pqt
SB4+XTMdd75/vbYwfT5ZpSwhbuq4UK9ULPh7ob82EenOwbZB3/J4q31vP+2pzEyFptXNVWkcW1c0
r0cLDdHV5tQcVheQBrScVDQs2dh7DaJ7ipdROCnNhrsXUFnyXS0FMZ4MY3MmkAXVdVzya+ud5p4G
l545OOcKfgc0tb7HH6cb9pITcEmrQRxRSESGhx9aKfYX6qS3+/qwpruJutGcaMEr9FG1Pd/edGMg
B+lk2zJV3RkhDCq3hJbIwItRxd/QUCcCQ4/UjydrvL2AYJ0x5axcEIRfZkfdU/6Rte7655FmDtb3
ZowBLCn23MPs72B6PkLROEeDlNYh9Hnbn1jHkiefcu26etetPORlcQfyU0+4iXo+Vlr1dRmuWg9F
AVhkRSNl8zbS9AmFQIeEEmK3oNSCBQJho/8QKCfN6r6ai/nYt/jD65UiZSKBJiOPXDcHRi3AhJMj
726GnVE4fhd7qN74aEgWuNmdOaWPCA450/qgzBritTzvzkW34OU1p6WE8u2izMHQJJQr+UboLhNe
lEA9HMA5UTT5E93/4SD6i31yFIdHVViArSwpGXUdFQucn1rTiUG6lqFCkmKw6uwVobjnz3dkYT59
TVTulzX0nlAef0CsEQ1fbeVMjqUQojIxASIsRimnMD9OttARDtYOC62stieBRGyKa7e9UdPAQsLN
7CxpXZP32DdaIXoLpCsV8QRroWzuqm1uDDdtONACMOzDGEdCG1+U84HWRfCIMEDGUf86oips/Lxl
xOk5t052fwaAi9dS2J8s3zrVDagxq+KpSXOMchport0SSve4GA2hG8BXz+Mi8LjorFHZBhQzRt7N
YpUkKT9MJGWv3gNS5jmxgee/pbuKBhW4mPH2RMowjqfw6iAujb3e4fRa0vhcGHBPIxB3LlTGCF81
MFW2Wpkgx4udCerC5kOmegKC186zw4s7A/UehpYo5c+nbDlEAhlZhwsGs/oyM7fdxgoRPIpjnquj
Eii5NSePB6JuM9TQPW0kxfMqvA2BdfPtm9acW0FC6boUKW8G/M1yK6GjaZHCeNBiVTwle5eWY9Ke
emB0PBtE+oJiM+n/hJ0c3lIZOhFuBo+MpKPknQ2U1BsseNiERjzcxJ5H6+GE476lPeSGbPkTTKAe
81O90gnYINTyYmw8moWpydXBNBphpinMINNhqU+t2FFCiDIdtV40P+U/CjSBnfzoulmjF8UrTGlQ
X8IZq2sV9cpHV98HQtDKLpcx+sVtWZsuv35YzWl5WA2SVpFRvtR8EAmSCbdrIvnt3bI6D6MXaTFB
3LKZFAEPRWim9TQ+aDFTfqvW2ZvdGyDdOX9t4KlFVPg52XldXKtEm+75wPJqlnXFC7jvuPiR6IhD
r2YRQpfOOl2kcurdxeEqZYcf9SudSMoz50nUfFySniiTwaLTVYLaEgB/YqUR2CP/e6eSo9NrA2M7
UGyO1kJGhew6/+wiurQewB/qH2Aj+rKAsFzrAPtPy1HR/e8Uv2QUrvzyXLmj0ZWLK8I7KKVrFBPs
agZPaanTLBm93aFw4Kl+unkcPU3Ez05MFDwKo8HSZ+Wchs3lz/w5Lu3OEQyVDE1KnIMsZvhh3z2D
mEe8LWZMfxXEafvfavRcRtGeqlFPAJCOobg867nhmL4KzwMjm938Fe01PEEyq8t2WDiDHKxCOVzF
bh5HTKRMR7rWjdGO1OLO2Tug0XaPrjebrFTINVQeQHGrjcolciu9CNf4ZR9SjhiAw0pS6LDiUz1X
H2X1tZyn5ZmAnMXJmhf82ukpGr4X0kX3YToR1AfxKwprtlKMuipuf22258mc1/usmNvTd9R9EHB+
FBUQeL0iuISIhZptCU6UTK0/d1Mu4v7CSj0Gi6wCF8puzEeoqVkq6dYPrHkXg7GgJKxC+m8DgSML
Pz6Id9E/wfmkFYlpFQ09u3lcNrdNCD+PZkBhQ4u51ArfWTGr7RxogND0xUow53um9B33HUmuQbBG
wW1hpG0x3vN/PjZDDkboa+8/7F7agPzUNVUJmHpbjgxCbUzLXBcMuwrAgb3KvhxwoFiQ4eSRKjQa
z8Q6UKsI6g9959pxNWw1yP+SUXI3tNpSNikZI50qkG0oBEjdKHaF170OO6J6xQ0dHLGEjMKT48Rc
ntPku4ZSW40T8PJ270O72OgAcKxt0zIfCyYpHh1A+EwOx/GK/zco0h7Xafa21KIYXt4JPFTM4OIR
PdkfbkR4P6XL4DMGTialtBl4ZumY5ODcgyY5TciZ9KJgzuEsAFeqbKtGEolkj5Mu8ULWiZiKVK8g
IuCMiacSgq8k3mvriyQDGHD2eMhUzvq1gXz9a1oY+XQO5SqcSvmbEOTwaRyVSOf2Z7ak68DVhCbG
ezlHDux4Rn2kixle2ApkO/en9avgFhB0APTdpHxaqu/UFIK8FEZErnt2Ae9d1MDRpI4XjQuJa9up
SMzPV0msCrzathpUF4AaNEBODr/lo/9O7ZxvQWI2BcBTa0V0podrFtNpW+vvZjSkzC6dDPVK/xwV
B2vVuZAmCuqAAPB/z8wM6MrfFqFojbAN0Vr63XIev41+U54/BpgavmjwDFP84P/MR41J/GWefR7n
CDB36Yhwj4tNmGQHXql61ky1vuEY9f7Hae/EQQIDxUL83znLYdFjDmfwpbl28ACjoXtzqbMd14Gt
kniW+/Terun8u+FH2jVaHoEFQjjrCU6cRHh0UPTaBAdedxVDrnTbEdzzEvbUH7dCV7NxMUmgcCB1
2bV16NWgx8EJXXHCwoFaDrzJYnYQPEDgILRt1kL6aPYjSJsv/rpuohGTIUiZw09utSysURnwpZdq
ks/S/EeHSroqu7vRjZNn3KFxwS/dPvrC0NY5vSxpalbO8H0gghZR2dNZlFbmdv6k3jBrccMz6udz
mu3xqMZt24BzuO8GVCqWS2JrpBg06Mo8CH3E5VKLUV701FGHGtJnD0XmZQhRGJJbK3RnnehimTgM
AOBqzzpllsFCAvxRcQH7kGBOenDhEJwyd/y1xnRRhaAYPTxr6/Bw4J0uJ0+PeKsC0DLHdnHFbbLI
X3/bNFQINiyMJ/h99s5T4s27CFE58NdGozkD/brlErulfDkFIoPnwCvWTuo6bwnA9V3wNi+fvjRq
Hv5lUec8fG5fyqMZ12OEzLD9kxDk9Ax2Wn/wg0bk/BNanKbLDNUeSuws7/vQHmTmVFbRbEtjEQX1
ywa4MrB+4CLdvM15XDUWwF7AjJ1oxEOtdkqYoQwZ6DvmNsrGnf8r2+1JAAqgwYqSJkBtYgqFPdux
JJ5Kf0CEmn/mlpFqcTe29D/i9T0LeT8CBveIUCV28xXSDRUqhHHyTTyzcgd8qucf3mXdllN2am4t
mRtu0BpyAfp5HucLDR4Bto1jxyV0CT1zq40g+FwQO41vIYY8vrCePuKzKHSTUi7cg/yEru+mwcMa
hIJHk8mZHSrnBZXXcLSViJFm1/uGJSjVYXpAcFPB6r0naBkHdwrtmW7TW7RbYr3dbF5/5aTlouWF
XN/7C3Phy7kdnv0wNFW9jlswivmh9K9PdUHnUnACDRgyM5mNSq1UtGmhpXGYPLcEfCHoKOdimlEZ
sfef4ce/Muyr7+a/5WgCI3Ze76kQvaAI8tKE3zpOjOkITPscFoST2O5bf1HGx0cCeyMW5qEm/WGq
F7bMMjnt2d/kcWpPLmYA0Ck9Jg9atWy4Y4q013njbOcct0g0tmpMO+qmAxMTLVrnERcHgxWQLFtW
rxThCr1Xis9yYI+Oir4CzRA7BhCfDLeWR34Qa0RThhCxBCH+swYqMEt9zgFHoL5Qqdq4K8mhuObW
NwNG0ouFnp3fidfPbMJ7EKFjv8ZaATtQ4O+IpnAti/gtXFimXLuPoN/0GNu6DxcL6ZGuKLGaCNQv
4IOXD+VJHaTutpHmykW8eK8r3Ww1L0OqjcI5Rci7vADHBUEU26Nk5w7wQRKzWY1OsZS2pBhCVU8o
5CIB+fnFKskjSczWbBWK9Djyf2xSaQEwmTRW9vgDXLkeQKdqEpWtQzNzH0X4eag/1mzcZ4ysKlIA
uy9dzBlQFqVfNY6L/LBgxtS7SdmvmvSgciCjWZyqPaztMyOUdzEdBm0DmzSlkDhpYPjocv2lBWjM
6d6wSyzHSWrmPltASMZqlSOeStMMNC5g0J+qawIWGhAVOI1qsaLhWcS8uUEdObjma0KPfkHRkZ+O
WIdU0rJijJ+F1NAnF3bJKw3sfA7OxMVj6937gMg2TxLFwU4GsN6svUcAj1i8bFnS31KDEQZYcSPj
cj3fkEU88usu+PIBoAwvSpavZ6XPO1c7Su47XRJWZdwb5SBvPKpvGFRuq+6VfTkwBt3PprJZuqZu
jPfbL9Ry/HwCzpbCU3x5Wi8XjhqpWfjG9Ro0J0D+7Sc/mIGUg3BtsfXLd/bNh/3M55wWABLDPhZZ
N/OZxb3QYDWYNTJ12dRH4FqHe2Ufu1/SyXJPWAIVwel4VbfVWpc/TYuJsro8umnxy20AAPymnw3t
zkY/AyRIgHk8sRCh4q3d20owOAiVX+oApvS5/YwDGfVduO+D7TkPQrJEy2K1cWCL+5YbM6LIPcek
0ukHibZDKrTWH2qUhOCeZoH97aLB/14z9XyoYQFCZHbCQI9fAfsrVus8Tsayk4QltLr5eduo/Mwv
gWbxNUYe70clSiCZ0zs3beKOP6+Zs1p0LTWZhz9/Cs2wkxAD9a42eaMIh5hCgkzYmmOmOYAnOVts
fHZzd8dJXPPeDUFIedr3U8PqFP/TZ2PefhGcJml4Ky48pGdper00JTxITEvDS7EVJzZX0cXfWEVO
9MOuFThv5VUcWWV48+8oUmJsq1Dh25NbIqPHaOzueh1izUTbRQnnhmMq7D4bNLb2VSAKkfR8B3QH
zzz+TmLXc21JRrQ7FaS49IzAC2F1u+q23l3LuqzkzZb8mxO0Vi9Y79j9Z/Hmb2lzun1uVvohuhFJ
qg+IyyBsqBkXnTXInGI54Qc1CQP0Tivl/dBuLH/mBRXtBBPiwyxI2dDJUkUgG98e3buRLJwc9QGc
dWTa+NM53G5QV1AORVnAFqoGo8yvpre/l7T3EGfvZ3a08PuCBOTB3RGcGNCydFcaRuEIlleXMMAa
o6ghN44v5jOERDdSDSzWkSXHIA/g6UTxLgBJa8YOw1TEQYZNBth2uHKDsyQfSrU/QmOd7TxCA3OX
DkK6N+0evHHvbaGa1SMpNLVDjsVNOp/wxYOwkkinFzf2uCjdAycJOWE9AtOgXSsrqtVislXDcQiW
RhDCIbMZ7H1AKI/URism82YCpfYf3xtXAMYNK0irZ6qzS2Azg8953Z4nE0WJJqbIY1hJdZxMsqRa
6tqpE+LeQdydR8SM5jjTlHIWAkC/zdG7TlIE4TG9ttI+T9L2qlHsO2gweDLRMxMp8BXkOoNdrR3k
JV3uRMDsSb6S2wS+rTPZ/ifNSj9aczbxnKHT43QdhTWAilssWmB5axjiIxCnu5lZ1UQ14o1YxBz9
nBA9mR4P0LmgIkAtqpkRQi/6AsGzffmT0l7CL3FFMqmmDp6HVVpA7B1ou/shvtf04qsOUl8Dbex2
j3TpAY1qqTppRIcvkitgLC6HfJlZFiR7feA7nxpJgh7g/5qa2nO53w/1xDofGTVT6Fj7swP53qWH
tNtb+6Gv+aQmuljb+6uWpfpmMpwCh6wDeymbD4zEgfKasJ1eRzdVr/nsbH+6gtkQuZYELj59GSwF
3r1pBAZ/EA8T3LtInAXNvhRnhEU3SsxtdCVc9RdsBlF/RJGK1WU9aagCXHIXF3nbu1pSXRMFLh3w
wP0gSPWUW+VTESAUOqQp5LUvr/x539daFOM4qIMXDJkWTwGb0p5wrkVF/i2JJM5VTpCgoKJpFODZ
caWn4ylhvVaVqRdnGsHN0D987V3mNUOVXkj5PEgw82Gv2O9m/p9c6jR9a/ctxY0/sND6ge8Y/jgk
dUU3yY2eQioFRUhSfA+Et42CJaJGMgP9al0SSUWcwtwZs93JrQNayNfD7Zq5fqy3ar6Wm9Xm4iCM
kpU3X36Q+eMMZVKTo7vzI8aNw1xvTWnnWZCA8m2YBKd5SPWg7/Ra1TKgcwQGYoeKn2Fml/3BcEaa
erlMspjPJ9CEJj9ypvvOOw1fD13fdvyVUyvaCfGkPZujRJF0xxO2KAUqSihMU5wE247UZK++ESCf
QXF5lD/wI8uim/smg97QFdgmtWY/zqkcet3vXDiX2g185e854MQODKPVt/nPtU1aDb3HSRoorz20
Zkwyv1gbLhcRKwWs4seF3G6nYqzCt3heazzwYh33bb01AuGNNzYhKKQLvibWH0/iR33c2/PdTcLt
gcpGWMyObRj0xGTu0t/KqK1q48rHzbyT+hehHpbNsD0/AOpOGP1Ushj73tHIBNtOy32FwDXx2jN3
6UL6kV6/QycAHMXBDn9Tz5E24cfBjvwoxvNp+iilcIIXgdDuUFxvSBOAQEOX++GSdm8NqaP/Z8eX
3y+h/1Q6MS+fnU4NcB43rQx6B6Q/zLbveMJCA9r1q2Cnk8NyKF1KsRnoajXpZXaCpRcpD6il6ni0
y19Xn/fDp3qx6AtX5Hfmtt99/uWSRUaIqiURz3CRgakl/Vz424ZrCN82+PdwFRWn6muH6fjVorFR
HSsTRkvtC/ULoOmnJGzfmz7ObTFXcGoppiLYQndMSeCoFnw4KUll5CBxucTm8LbSLyt5ELK7fhLb
kT6svgyKzRch6HYvWMe+VAHq9L7hmZAQ48Ej8EGUYuIALoY7C6zSRWCgeIKZzOtQb1pF6OXc1xsx
CAWiIkuIAPWOtOPAbH65Bj2XDAAN2WdKz4dlfSi40iMHbEeUcbw4Km/EllCNYkqL2Iac41KXx6qa
Yhd6gENN1CPPmBPcvx1x8fnIQmoai9T2Qx6w/8UU8WcPNHechE8+cX08WLTdQhARklBVsbEUyFqZ
Dmvra4dMyV1IQx0/U7Bt7w2O0k3iM/U8iJytz3AsQaA56xD7WuN8zq6JnaY7YIwQeiufsHU3Agpp
dlpSGLO6VPNsuXqDVmwRwcs6mYwyMbtPIsAd+JS7iQC8XFZEX+yVBx2hxtjS+UfHO6QH2kdzgb3a
32SJlz4XS4IwKP7thCwfAgPLdzv0O1RRIxzaa8Qw7TxHeBlVXhs9L/y8fubHeEMxUuUKtxPxbWhH
tN0HJze8bJWAfbyn9HKyJlzAupQOBrt36g9uVEMyVNeOh0WIsvVEdM5a8oU2VGamFoDNpJOd9ywa
OVj0AHT1CoEuWHIot9tKzd9Y6ssxaRu/4JWetgbvbXmS+JsnDRYT8MHSJbo7cNCS5Q0hwCNrxUt7
/jUeMywpXvW7722rZQPq+88VnKJNnmg2YDnYe57QRP05g6VTV3dJyoXeYt4Rl+T+cG8Bk66VelgS
CZtTqEb95R79cY0asjgLV8K9VDI1J3VnABUfhyQHB3uO6pE4IICqdAVSre3OAl4rfDEtra0rarKw
0RTtySLVe/P8VPnE/u4VG78a28AYZ1WdS6Jb5f5BdmMSc+lMrD+2+9y7C6fOw9vQl2iefGVHuZ8A
KqzuCVvzXm9LTyZGvQFhZW6MhDhQuEKErtcfXhVRBUwQ2I5Rgfaz+QEjVhWEWhRLk+/ab+yJffUb
58twmn7AvHUYFVB22oV2yYuxyvmA+nQDXWCvLO8y8JIvSppjNVBKkFdSzVpLoo3gLuNAvqdNIhW6
SUH0H/3C18rSqbTybCED1bnZ8GFdnAZ9GymREEtx7yrZfcYYN16zIZyIL00aEKAUmwORPa7CRnIL
HJzD01QmtvDqgMrbRl+4Lb5cjsXrn39/G3gWjZ4PKdT5LZC5ETqdF19BxtDVMXmtv9jFc3RbIdXW
yt7Sj7Bhw5K2ACyPcOYg2meU6+inLR89IEM2D6t4ly6sRrqEtEiXjzQbYzo2l46QzfdMgErQ5jJ7
O4S9RJPVLKOPbab3vLLhZ2OCWSI/TBysp6hJnJ3ecAy70PGQ9yIG08ZU8E6gBkvzSRuEIxPW+vSq
oUgn4B1ZetRnr0DOB9sL7NXX5QdMrbUpmQaAlmHa6TgekhzZimxIC2QmpninNDuFZKhSuGB0vJE9
djXNFGH4TSgJP+2j6ZiD1KUrIGVhzYuBt6lynmqeFxVeus+/HJTiy6W7AGP9KxbdNuCIx0SRJ11c
UFGITpNke7skFtONeNN3ym7A5kT0d+02N4Z8b3vaz5w9pOpH0fb2Qk/1mOiDjuElxaciXqTf5Cjr
IE0Rc+hkvecb1LJyqm3/3fXnUfFFAqWhCegat4tw8UYuLGI13GMe4Myf5a7MGvUu9E3eXqL0zJZn
+rzcOYCPxGhfQWwODtpXWuCIE9IUlWZ4MAOmZ8VbdDwUCN54qdfDu2oseUe+ADS1ISuaWLKTBzhv
gqjqhVlINX5o4+oEjQdfD22KfND/49CbR78l5iilL5ux25mIakfJKhSlmX1u+abtrL0dVt/ClAa4
m+aMzyF/MWW/YcxHwSsKNX1iL/rjftjKuVZDWVpnBEQi0fbfWzg+U+SJ7+zE3ZoueK1UqR4vw8tw
YbTNW9J9E/7WJxEsc3myWLePHrSXrkxWExMpUtjmg45Z3u1FI0YyRt9bpFXyNYS+gRnujBA/XdHp
Grjx7MM4/Yjs32HJ7E9rzzeJVd21WtJ+asg5HxuhRSZI1aLsj+RF/IUnvzQjtvVY8boq4jBq145L
o+1qEWV2mCIuJhgz8eP1KSXD7BrjW0ljTFxkiZMDFyEpvNOqLIgkcSQPi19Z0E8Q3LqWj1VfhVLx
AZV4uk9gZF9IQ5vOA4GqXfrYcfcun8AInWNIkTKVrVN6zhlkc1K/LJzkCqksALRXbDA8LCpIq/w1
KKEnvy9ORZ5j24E/CrODhdG3vO7LRTd805WRLH+5qnfD8c2fG+2g0B+EcA0m55/C7OmzK4QoMq76
rlnSgztI8b1dpmyWCrVw+1DL8Hp3dWCaH9CDHlPC+KaOOJJOCcuSrYERTMeHM9PRoyyUsJ2RWArO
TUlreNz05qeteyMxqkE+CjN3+T5xHqn4Ie1kkMD6le/UfqzCZ4My/GcqJIt7rEbNISM3QFusXBWO
lPK2XA/8wUYDSzEVtf/LiDLKKN0M403Hjp2lA7m8IRv0QySLmh6BTzBNQb7ocbdAamNl3EEFRwTP
4mOtAO32bBU+hNEMNwMyi7iqLbMALbaWayCJe9d1gEbl2r+8cG83AWvYbHhGM9PchhvuhyGGQqwn
RwHXEndpYdTcMjYKoFIomVB2B+hsnx4Uyq+0bZwzW1ipVoUCYF1+R6ukAtFfkBs30LbMldlU3PnH
NpYdiLXt8T6ITq99Y6mLAGlX8CNCBzKVC8RmU+K3AWsazUc9rw7nev3FSLl9w13oCV2NAv41AixR
gSlLGuQRphaO+f75PaSJ7P42K5wNEYK7R+rM5SMvyGmo34Gp8+eEwwzzuuRVpiQ6Uf8oPsXICS8K
ZpDDLPuU/tyBhEas140Cj0Huk6MTuveMRJi7QENLwh3mbIpjO6sRR9qGviR0kLXhSPMWPpkxjwly
3Rxbol1fJxHqyBIiJlgiO3FoRwp+Q8O1/+YqtcXMftBrSJGKfk2j2tW3qIN6qQhzFbvoKnBgzI38
ePA8396P+eQjeofcaE9zs4/zZQB/bQrFSxT9vkKKF/aNL3MohbVzTRxbhdOoApo+Dwqb9GFSZ1wP
kMQUrd0F+nicVVOpFi0N5HD8kyWCGp2QUR0IxZ1/ZXQ8BzgdbmE1+VAHggZHdp0s7ojhNty4ZwrR
BFA8KLlwdH+kDqX8AXOlfTjGDWABTEHpot7PQJ6gv5Or7aNjJDbPT+x8wVxpYp/tKAltFRl7knrU
MAuboX2x1dYZJ98SOeCd1xa75H6BX5j9+4Hj9w4GKdC6jYALH84n54KG0QkUMbEqZ9NYj56UWaSN
6hm3BQJxupFF2nTO2vL1tGnkj3xJBoHSlI44kLAJel+egFpRdBMa76ZVd4ecesYky0gleqdNJkfO
m1YUprVfsWqh8Jqd04IRKp41u4k5dDQBFGu1mPaZNVh+Xlq/xi4KKKNDk4+x2aDIY0lHnd4mzawj
PPKiVQprCkeIwpwyx3gImSMdgzjpanJSahFp4CNZXU8i/8rIHqhvN4nAqng7ZtuWp6JbH1ilP2xN
+T8ZQes20+fgZGugUaQRMtrJrgpgu/BdqF6K44/L9ZQpRn+7Caaij89U1notcAE+G5BQRF/ACOAz
C6JiTd/pa1NkHfv7PNLhJadVdr4nD8WXyeZ8jNt5FLlITpSRzX1fZV08Emmb30O2qKfDQOi62zXZ
kO2ISdhn9mC0MuzBYkr7wMueNwIxhqzgJD7a6mvUiGHP3OLgM2qtkXSJ1WwsDDoQeky8lznuEx2B
N3BiY8JjokY2d9hXAsK4fNN7uaQib0xVMRAG1KWpxXe7miPoVtxxm7FSuM2HkPh8L+eUJ7lXwS4a
k0QsU49TDlkFk78eeQpPWLEP4WHV4q06AOA8BVna4iSlCq7bgtm2VfzsbLHoXSCsCveRMZq/Na0i
wTN9rXLQgyf7br3ZxamBF3mV9+Nts7qnj9JiV2UZ3gz5v6Qesnf3fpWAfb6bWxtljb0WTvguZZFf
zDPhgZ7FC54Wf07bxUR8NWm9xPYYIVjSVncM/4LjMbSt9JwcZFLazHvE/CjxiH1SSPlcon8dNfml
1GWmnMBmcOxPVP/T42RB7MTCaB8us1NJXVVEz7lZMCwyz8DiDKWtxToxlWkiRwHRcnbEZQlRydLp
LNn7O6lLfFh88ycOIUZdTqt83uR9DiMbzjClcPDKS9pSSOy/8HcuA9c1l7Jp7XYRftdupu6ZEalt
Gxni9XcOAaE+niqtGimfU+VUxtH5zSK4Zej7onmYAGZsPR9PS7GD0XJvh33BSCviOzn7F/Vn4qfy
pavUyA9NoGRjxQkJXT4J9wfmCA/ytjZO43ti6YEAl8I7xO5zgql0Aldbh8JrOwRR6HcNxukYghsW
Uivk7856j6XeL0Ohnf2LlKFUKXOZu7BZN8pt9wgsJrxB8eEwNPQkA3U4dCvuGjNs6RsueBZjtHsW
zrQYw2lUwUsxW4Yt5TqToBwmcXhXDj2+SjuSto6Arg95goS8EvxIsQfij0mF2foZfrG307/N4Ks1
khHCAaPaJ3A8+WG41kdoFxal7zrnn6+8foG05NY8yPZQOXr5D4Um4wd802yygjoJFL+kclpV4Jrv
/YKP4JxbrsOCNavrfEfse/quNmVXd9o2IBB7kLkXkWYzbBsrDk7t38uD26dl+gTd+GChRaFNIDK+
A5PFDaprWe/11+fCKzZ7+vb4PfRJvviz2qzUHGq6wZYyy6OaCziMcOvk9oMZWi04oEgL5kkc86so
U3Bgwtt55yWQp5wheGypBJjKVxQKyd+5VLsEo1pTZXuSzLTTdP4kDlAI9pOeEh7SYggmQhaFPNaE
uomxfq0iRDmFfYVGyMFfBwrDrjMGvluwuP5ShubZCUXtvXlHnjrCZcSlb6yok1x+LMscS7F1Mhux
OHMaerJ2br7TEXKQHqMdM56vDXvLTaTDDcocFG9vC6N8gXqug6yHCN0TY0qIrpY8aRioYAm2nm65
ojtjjYDMOuk0Pbkv7m7d73bjWcaJqa8wNn6BuJfCxX1zEcZLkGupdVq4s4IhLYnnaY4YuaQcxBWR
J39jq2Iw4Eq7eoa2yRRXYrGgNOn4gmtI5fH0di/5mTffuM8XtqnEbeJTimMU673jxEEXwTYWMc2+
UxmNC46sYf6QBsZoWDvH2T2mf4kMiydZnuJsGftoFSlzTr4bc8hMeVKGfRy1VcPsNcbGTHHD6wxd
nfe5F+ndfF86BhS2ese50xkPFd0HmbYMCMWEb3miEGH0Ntv4DQHNVwmodKefNS9VSv/jKfWC/7MZ
swy+oirHSUj99f9qLEqzIT2xQa2Gwxn1e1vmJMqfrm3tLP7MTBghMQYs4wtma9PBYut+7e1fPo8M
mxKkQTFoSVzqcMYxC25lO8Zjn/bIX+raNrzCIXPtIiOQqOBWlNvcXs1Z5AcJU+XRlQdoi2sYWGIA
Xlo6KaKy/56dh7RUl4xD4um7e9UWq+Gp8N8Sy4L6d13n12XoQ4DrzW1Qo086buEW4AW0JlT1JpZK
d1T6CeSIHJYfJ+rlQMiWHPTrU7VHO2OEHv4BMVuhAoVMmwU957hSq9veo451gKvtj7IyYWTpkKuW
rGb1RgPkUY8HF4xvcVS/v1CLITopT45qiv/Ap+WIn8dTFbXQDZkD+pBWoMH8g6GbFRCU6a0LoswA
dgPrbsHr2FQnuFiZHvD74ufKA/sbEIzGo4KrrgEvDICX2wQfN3HhBjvP7FSlqmVRySzzULYGEl8U
nWCjSa4ZFxcy7H98GlWWAs39XmCOIjnz15U7PV60rJvmoAVT5Q1Shy7ZwC/ePYaLtKgRYdRFw9w3
QAoi+CFCW3624/uT1x+/3AOgT6l10wPIyiclN/jmA+htAYWoJkKCrjYaSw64WEq1Kbg1kdUm//L4
DuOJUsA/uXUu5L6kR8SQR8QJglTa5MYnJZ0hsRXGauuU21WsCxI8FMevawrZCQydoQIXpT3ZTr59
Sg4YVQcBnImnT9KT9chJch4wb78qZiJ/aXb6QY+JSd2qx8PnQGax7BQzzj6TZnYixYNTPD361W8n
Tcd82Ian/4LwniH1sLRbbOEITTDSTDkSUgvIOvYTFxqa9cxWtr+0UGVsrVuuuzo0lWWlIygaj9ga
EBMfd3ZPgSGRBH61n95kfYTOpQKg8RxIyLXdUIHpQnWLVgpkqzoCimdbRwR04PElaSzDk6zfx2q3
xfEIuXveQm/JHKHmFh0qJgdKZI40o9nlcVfN6crIMXoiRJhCsYFK8FS71hMdiquBAmTsLE3YoXkB
XhWPRmp8hqxyMoWndl+HZ5air/sFLGgf7ZXrZ7rj69u4i2RRudtR3XKcmWGA6sC40wCZSmO4tYV7
R6arLDGh3Bt/O5kCKt/xZQr/UO4U5cvkylnMBu7l/QvrcJha7L6PR9wEmbtpv3m0zD/78pX4dx5l
KvYWGYvqwjjUs3H9OCNUZ9fd6ycQQ1V6fx51d9GThAH3lCVzXC5M5WAmXVidSJBMQox1JPPRr6Zt
1tvBbKXpY6Uz0m7vwPz9Tz8JgkQTCCwaWSkp07TEUYy17Jwdc34H8ty8jhQ/ok3mC80SQgww0myI
eQi9gBCzftRe3TshAI9pR48KKSX3r+bEGbfWgAuswUp9ElEi5SgmFCA96hy0CoB9PgdRf0cS/7E0
ZBtxkGmmkjNOfE9SMfs8c01wdZ7nyVxazpXrlu+SoM8LiCZjR/tAs4tJpOnNqIbG3Hv08DPHv5tl
l+TlkXwDme6LRDpmfk8sVMNT1kEAJjq1nXgjWtHjj4+1EyKx4W0LtP9xlDhK1Rh+C3cp4ii0o35h
CPStFdtXPwPSP84WEqzdYThSQfdQqiqG3JTV7HvrrAfe2sQuguKq2Cx+l20f0m6D2Ok7zNkr84XT
DE6IweUKFRgqZJ4gG/CtOnDyNTcqCI8jQ8bsYE/ypsTj9kCuSqXPzVB6bbqtp8ImjK8k2M6GIWl+
+dVQOvU2n5/LMb0wy+rbkjOIRjYSnPV0Z00SqV3gZibidrpx04NUz29hMOJr+CWndZ0OxOGLI8TA
UY7C+mOfpEuLkBIiUOqOx2Q6g9RXKdljUERBaN/gXFfWTrUQVjEaTiVb0NRWXMNZCeCAv5DVy1Ut
gxiDvZ1myOLfEaB65DXKPhOXD47xf+9IYfDOJoDG+kOUjjoB9GC297pe5GdDYb9cDmZ06SKGOKRN
m3kWm7t/veilewD42LFhrp4hczugyDirC7fXmSGpVm+aN9j+eihwyD4m720YDQgZaA5q9r3T4UZZ
RH5Jasjc1WsqJ2PJ7djZ4iRNRZHoFeSeo9q9PoYpC1/aeXs2yYm9Ls7I00A34j82B/Z2tBnFoV3s
XICXDG7qP7pAftHm4m6OUfMBwtM/zNoBvlyJV2kmVg26mMTdmTml05MIsrdyavEuuhxUWBndqYAs
pmdGa9DE2P+COBPEzl0hs3NyKu/Z9Z2+yx6T39HHtRz+v4+C4bTrPI/eX0cFGpIspnNFh5xpYPHe
8b1gAT3ekLbXWFDQagXYs14hwr82KZHY1zVka2KHubBaoQj9ToZ73JWzJYN1SV91N4qqHWbfha3b
kutpekyNM/xRrTUjuXCkYS52QRx1FQrgYzjQX7odPwk8inIdvLdQzd/PA9VVqGmwBnkn3rhGtqzH
k2ATNlDh/sSYIv0ISztYGmFbopGc2Gs8zqNAPQLV64yj+ZjCLJu8K4L/2vv3FbqYST66n30wcLmJ
lwx/Zy+HQEDORbbwtCRYT2GS4iWgqgqC/JjEw+yZI2K1hEWRsVJTvIbMiT7nlwbSMDf80BmMUeMx
Wpa7pjP+woJroUPz/WD6rV2t2XWVcdVr3h4eLKNG8T6G5bZ7Bfn3ovb+FZQpaox8NBh1rVOjZEGT
04sOtIdD6DV6ZUgzxsT6LsgcS8IaWFMDFTTjF8zEoi8g8zrcqHcOcrjS2FxaUJoJdi8tp7y7vM6H
CHC9n5KZ8VT5zFM9hpt2rBnXiNbwv0IlERxiNqmG9x5ww1iX43TYYULPVT5PFOozjO+gHrXIAfTA
Cjrk0eKnlEWCrIbycELWYhfUlmtMSRwndygl8gvMoUh13gaZStC+n8HAR7f/l9AKHY6YQu90XdDp
8kCaeLplQHj9cUqhwmyxAv+o4uNe4Yt9/HFjqhqCZWXH3E0jIa6WzPr1aL1MpMtjwLCkJfV+DTok
2gSL7Sad9k93VN1BSE8UQ4R1GWToKchXf6tUnjc3oUloD7WfOPVB0onAEou+RxzLoywPvcJWI6tq
QEllgCLjFXKIJDPLY++2L4SFKyOc74iMFliZ5gKp2OqEYLQFwa6YKstB/vZ05Uggm3AHFhmDsC99
412WVSr/pK7ChgL4qWBd9BsEXqApDlKwe7X+vW113UZtVQTT9KESzf1Yd+6lm/p9Hjd7hBtvwuhh
V8ML4Q3gIdQh1FM4VQ9vm2/lR+rA13wavH2B252fSiVEpaKm9g6wJbPnOhdnYHPXtecLfj4aqfDN
hryIRP3HXAg/T3Xf5T+cpvsY4Yx7jFKUE5Ap+tPpiGoQApb4WCuiVsv2aLF8R6Rka8saoVMDjxJb
kq7zTqyKOLB52PHmREMv47r/gwCi1VANhmhkiVvs6wlADNhepMv3du/80yAFW+OKJK2oy12/+2Ye
nSwPc6mzJyTYdwmJCGxU6ClFDIaBHUfP/8bdfDdVvVIlF+vmlfJE9+UtOqZgrpnPfDw3NbjaWl5q
sHoj8HDpPGfjc+T8CdEIMofcDmCnJScKLyuXv2MtFiirnfZs6xgG3Q40FnaFe7vN1BvVzny/jGWC
zh9PrVRTf5G8u2FqWr+VbZZaSE1r+R+l5tyfcfTJfni3To6wK9h++UH+nmVwYlxH7DFznCzsm0fx
9A0pWc2k/wS+V6cMHOzsXlxDlTb4RVgQgbd9EFVE0HJVXDlDuQrR8+N3Cd2fHvaXUMr8Ge3I/EOf
3NL2jsWl4MnWbIwJ6GEIOpqs1CnjNbdkLfYh9ILUgYzjcwsSLfzNx4aL920vNwuNDVrVTuOSJ7xo
1bhsHQ4t2ZvfVAt1QV1vLFzFsJMtytSPGL4gXoKNeBbO9K5etVkPG/gKf2cpkTNCg6a+g7erh3xT
HL49uSEFTMdHRxOABqffJs9EwmFIXTHOFpWqbqBcs7ZYiT+Qcbxig8YLOB4+1nHYH5dcOjoD1e2H
boW2BPP+12rc0JydM7AchLfTG5pQoh7ie/8VBoMFPyFiF1DZJO5/wstBwc0sXfRGv8BKlnwG68ma
+4g5+nwCpY7DkLJcSYffxFDmOfnzeJVoLcALqMXYEcDaVOH04cnCF/sQzMrpd9BxSwtYABw7Dj+2
Fj/vOeeA6hv9vTiq1Ww3LSQM1vL24+hNB8q2eRKdu01ZInhz5Srm7+u/5Qp45F9K7F1vgPxXrA1/
bg7jKTTQRzUX4dPKIFAW1j0y7JhU4miEVzDQMfy54abW+UhS8TR/z68E0LLXoaRL913s/CpNXTvA
r6XeW4V9dSuRUUZH3tKNPpoy6RVcoryw0Jq7dm3AY4rAJT/b1HSyNCICfl5n7uFz9BdmTofOqYcP
7uFe5nwVSh7F3GAge+NoVNW7UyTqFy/9pkqBQRBfbUT433nh6Q4yM6hPEskFjCVTWtVyjXdnpJK8
VUnXj6szjFiwSqXpUGKEbMfKRALJffRtMNLz84tHXSZ7O8pSu20flXXF6dsxmrmvt7NYGzVyEQcV
iNuReNKEoOxkKL6eR4xFfOmDOjD7Ibt3cJQlI+KFOCpBKXCuOmyhf7CS21ZovsL8TwpqFK58cnXS
253lN2xI0Ig4zW85ynm/kO4e0yVGrVCHZQscU54L0GTjf3QoFcLNF6cPA/5OzJuttctaW7pJyQnW
Q5cjHXQMUflGHKEakITeFV2BappksD/TdNfRip7TZXXW7dR4WKMXp59K8h0G0Knnpku18k+I4un1
WGfqoXhbmVfFax8LC06rBQ6jaIxxewmRwjgIVxiCqP5gsuppxs9ujJSqZsmDl2bQVtKFCPb+bXlJ
Jk5R0+2e6PAGIRLdfu3FLSoysRH0WOEyW5GdaW1urk8gbNASYYWZCLmkXUP6sjdQpi3jwdDP7xaG
uLjJMdenyZV4N70V35qL+LlSjcMqycbW22uZm6xONFV/SkqK2NZhhQCALZIaVLsJ3Yyb7RkNxcmk
RGfZPS/GKAhok2OgPrLMs5unjb0GNj1JDklRK0FwVFEsoxby9jkPj+UApvX7dlMJ1dNHEhN5Krfm
m+E9zRbZ1YWGj+iO0j3VpC5g+8CLTtrD2TTLa9amFi2Zkr8W7Ox9E50UbXxaQpTjpZ2Qy65Rf6x8
t4krD/o0YU1rwV9mCt/PZFIeb2d+kt36fMsDnDPjK4+L3RmZocrjOhuzXtyKTUh+494eqtVPzwyF
zLp4Xsmt9BZ5dcPK90LNtsj7n/HDfgU9zA+q8TPMRT6bzDvAoB7yDiE3CT9dU3AhFflRtI58Zxnw
ph2iiQWZ15kjFZZteVTphreCrqsaX1NAQ3HficsID5TEZYLixw4P3WBSHkl5cqHU/FVw7qP+7HSC
hxG8joMTYMxWqJcN5HE4AO/RH+WcjXj8NCSnIwE6JOssG9SUZfpZnXJ8wENjl8bbCwAyfkbLZI8E
8OT+tKuX/EWaY7obJps/jOvOsTl0MboFK38HKOfBbDop7mXnUxuKEq984Bx0SWHiHsb9oxrFGKfo
ZzzJ72eyq3YRG0ClT3EXmpfVmPj9ZZBC+gvpCZT7XhBHGkaSAj2q9RH9bwXtI3OfvmRaei7KG26K
kI+Lo8VMuPdsnoyA8XKwsrDebWWfPX53U7d/R1174ee7SPxJ/G/XhwENIamwDziHBUKHxbVVq5zD
FxhoMQZEU9HGz+o+g4tFbWCKIwviAOwa6UFMmZTJCF7JqUwnAh1FV3+SX0/4sLBj8kRe9BB5i2sN
UvHjy06SXvN8ymM+IklfTsm+ccfhjkzq2yKN0DMKxdHuPFjy4RzT9R4zAK/F0ohpl+x3EZnuzsuz
0ots0cil/7tOHHiKsLtjpuAL0nKPphCvbRuiEpVe5NI4uNvoYRigIsFXDqmpkGGyd0eBEgPbcjAQ
gIIHTYiJ0D7+mglXNv6TtbNHRMa9Axi6o+HoQ4H6J+8wt/+aaVn8l9Y/UWsUvSCmFY2y3Hfc5zJF
INqI23SNMP5oawTSj1wQoFTGhppX25Pz+3WebPZfEJ6CTxdTTR0DHBs9lc5ZcpXCNKnTP3vWRcri
zCKaM+qHAx5zngbcPpv16439PJPxDNYu1XaihhFpGy8WXkQ6Q03gJ4R6Bhj4aVPGlUX+umddYIP/
YPUeIyJf/CNsVlJXuZsWxntIZe6UJBexKpHlTpVLkrs9rfLaPf0GXnD7XXu/G5xNixjqhTAcntNa
avT7ws9cqjIwve//hQqszM2I2M5awR2xjeZalxSkvYr9x6VnzyfaJV9ZukqM2c7IvxK7b9h/5Y0q
FtxPkaLwLfYQGXSWS7iNzg+OyG97hg4MCXKrMsUX6SFLSzIsDXYbpopGaeum7VdSWE5J3aRRNZXQ
MOG5zvvful5UOfKCWtVGnaBnF8uGzOh8Vnb/U+3MsK6YiaNtG+Eae+fLpSUUV+i1HhdDV+4AvBd1
ld634ZZzxxtIubZtLTWXieM9pgoZje+5CPjE3tw4yUEvO5wfhX4J6KxtV/C8a+R9h6Zgv0nCuJjC
HuHdl8uP5Nr8f/28N5zFtC33RfFOHb4g0zZ3LlvgFDUMcw9x6o5q66l7VWg6Jo5J6GwaI2oFTGUH
aKNlyfEeNZcFDpQGqt0qAlHAe0fxtDI3k9fWuIJaeQZoZjTXHQAOhmVlcLtlw7AG7AGHHQIz8q4a
4eP3AqamoloAUl6Wz41jzRplQ9jLWHanfLv5Q1mDiGpOBxnNxC7Y64M8V7zWzbxi7XXOhwm+cQcI
IrEFs26PnXCZDW7NCf9F4zfvNfbKcKqofYEGeLyimzvUuQoe0cXXQnHkA0XspWd4uOda4LdyGsSR
M1wDgydYGrplKFzsrL1WJHSzTN9AjkfQJo7CDbHBNnBXasAtjOXhNYP5+z8Okk8nP2RUsQK8sATX
78M8kDmdtGCkEviCC7WQiUekV1llo8vjAw2psX5kUwnlLShNsqMiPQOcZEonR4C/Vxv1Nhqx6NfC
BPTd7Dpp+LnanvzNkSiJoa6VUWY2kFpbM+GO2vAjCnW6UQqZR9ztmt1iq0Y1Jf7E1R1rYEKL23l0
W9tcNyZWGNx9H4Idv1cZ0wADQ8a23jx+q4Qux10ZlJcMawPOOjKNihc48PQDUFn6vrgqw9fMsx0D
HGEJzUrnbrmxn50hK7cPijyVcMZnOBt6VnELR+pbhOACIksVHqlY9lATKArg6JVhmN4O4EyoIv8I
kFZre/4gCdALaAu1UONn9GJ+OB4WlGXi49oFcS5hQzvUL0G7UmaXrz82QwwnOklEXu+n39fFN749
FujpIvTT5ta2BUmuPH0dU+0GAmIr9PaghHMNckieaoRCAP0alP9wzfBh4yrdovf5qLHHb2ecHzIS
xLKTC5AMaYF6jWmWhtVmRN4fe+NAbQk5jaMpaVutnizhcy6mmQsKcV++4ECsuiEI4JsEFHwmrTIS
TDS4mKlo+8Gij8FajZls3mY4DSkIRvPGaUAYWl+k5Qm9q0Rw0BRFMDFz7Mmk7SOiheHe2c4g9fx/
O5VVpzmSZ+OW64T7tDA9K/rXAl2pOcdCK8PDPWTJfTVud3XM6ufAhLrElKL5y52QpLWZ47Sv963r
OUVjZkQmgz7cTUXD9f20Ey/Tkaj5Nn5P63fzBX0FK9ePLPfodHjFsupdtcgOfxUzJpUGj4qba6I5
Q0Lzy6r+S2l1xkVLNo+zlzYk8PZ9f6XT3NQFpsBhLOMiLCOdds4URj99wKKORrIkc3F+YMgoBVkA
cDxKcgmb6ViF+9FKeriybD5Fz31YGsKR06xkbOar3/ouQUoEJID0ERw3FWqeGr+uYFfuVJvLee2f
gLdaap022BYY4IAj0hadKS6fcFsN8abqsVnD1k3xbJI/59sDjFFXNzKL0bzjhBawgBL4gtec6rW0
3NjxMK+PSCslf93netG5z8+6vHdVCl275PU7bnbp7mcOHUlQ2ertJhbgw1SL7b6nBGVCPE7qX1zw
mw7uuiU3/cLvfzBpu9qimPAj7ue1INhS6URldAfE2ZYNqNdiOsvq6u/Q2ulgdzIw7XjCd6GyYl6I
J1r4xSPSIjU1e+5zHKkVyvw2dgTecIvVy7asSeZs4395gAPJ3PjySa3hDticbtfD4eWKgsrp9oHp
7HYGRwk1iDWIhf0PiU9HES+i+enxyzk+lzB+ldfZKaT96ww5OXl+JK4cJ3XJBk4xTnNO0KIgDXIe
RLopDQ+R3URZ1AKd2UScAPU7vBVKIyLOQiVRJlWg/eNXBfP/MIoe7oxkn0nPSQkGqdQ0aZufwJHL
xSZsxtkhME1famUINblA4BRkVr9EI1CGkE+dYmLOxBtaKr9YZinsPtlHpPfCmtHvAnEdhD+JPyau
q8+a8btxOJQrrC41OCFTaGyi7gEiws/VS6crucyxfaWiJuVxeYyPeyNpoG1+U+PlKPhhKDVALGZB
49AU54+bJXtL1WITpyazmD3slVs1NjbxN4ky+hz97AFTeRMO1jbNc3pMlQp/dLsh4rAAX/fztiZM
VzzMIPagqsVKLEBIaHdTVcBeKOxMl2QIe9AHqH2FArwE27kRcY+jWlKbyvYhGDJBqIsMuqGGQnPj
7z6wEel88iQV5JuoFxCjpTP8Q+l+Aon0C80YtB9n/vTktlbqAnjux+EBNjOPPZzwcQCp886tmzNf
xV5xLIVne1ovRISaoUE4bRrRkslivSaTt95/9Ft0qWxZvt5Vwe+0pU6Q5rzZV2UpsybMmzvwBBB+
PW4rkMpJOIOriaEkfObG/2DhRSQ8FNabVpUrIiwj3p61AVspa9kdVgomVvLlpWeC1IDZnbd7/BGY
qe900EShf5zk2xSgyTyoTYHS1jXp7BIBCxYiA5Mo9h1hx/+ExE1kR+zcRvEhM6gLWWoN3omoQroZ
uiBvOXrZwYGohIrwmR7Enq5QtzbjZgcjwZyR7s6euTxeNu/KUAHpRpRciKN5Uvg1yMLK8RIdeQJf
CmFWacR5s9YHViSb6AoTEfgoqmdOm4ZwFz0FpVOuxnOIQpUvNvbiw4s/1Km0xAqKFmwaqx1Z0Sbs
IzyFqPz0q+DbsVBcHplAIK109hvqvsnzjRkD9tkOwV3dGGvLbQ1OWtHi1bMbBB1iuSPxwDASjG8I
wt3a3YuPz9P+9DWV/TYvtgHv6Q+RFRsFHBHspfmGSm+K7Ar7R3XSuZYBr6On1i7FVEDMF54H7rV9
+mOW51AArDD+wN/0NVzb0Mx94MAqxvGU+gIgEHNCj0lmYhaaeewdeRVFpelF96MvUytgJyYz8Gw+
HpjkhttT5QkcLxXvGM5QG4b1o1C9b8yEES4r9jASgGiBh8ptN12l9AOh+TGKOxNXkq7HQJDRca1x
Hp/Bu+mfkq2fQTrVUUIz0S7tHK+UfV+YoVhyGlV27S+070YPS0Mq7MOnOCXjrlt6oKVx/TnUAZN0
lsKUSSeAE7hy2pUtfQk38PyTMuLs6Ye5yCYwfsUr9EFoCi24T4OKyrE/lQP73uhwpltmWdsJuvCP
W4udTMQK/0Vd/UOXHzIUGhPsfGES9YvGqm+8wUJ0iejQlYiG1CtM4kR2mn1sZ6i6Dhl0Jby0hm87
gs9rs2Me/RSf6Pu8lTBjEWutyiCY6+klzHBPHw8JmuQJR1EvWvmfBg0QO5PXiu1Npitp15CQOHGF
isxeEuCijAaoNGkvZzWIhQuXolbc1PLxIxJGvixfBWWvg57AcDwuH9tUfE3v3D7wApEuUzgkqV//
hYaPMVzv0Fe1dt3QydpI+SKAJ6a8gIky1MUZPiLVsfFYRmZcdl5TS6FFWuCqeJ/oM48G94Cmo0cE
gxv1K3HvC32zHqJGYGzvd9HqqDbOyBhKtt4ErOmuHPN1gOZuQZdq979tFY9pCfyeMOvrN/R6i+uf
mArNCdi7ranDeuM2tH1ocIfRBgOsNvKVbYVD9XdTuLyj8w2Vb3EiN6qYw69KHOPPZlV0iC9ISVhj
JZOqXCRHhBVsi46YOw0nCqCuH39TDmhnnsVDyISguvDrFaXwdwpFQ5uRfBQBHO1sva048weGMCCW
kEYPmboX9lBgo5/2jA5pripB5s2aoWp++NugKyEdJGybGop5C6tdQYjM9rkgzOwqYOchU+k02iad
mPcFUNKFHZdtWDSldPrEeaGXzyd9eoJl9R4Kj1RczjSArZ+9gBmRp8VMenOoZRmXjLM9gJXmI4Ct
OVKVeLK4FAitduMgdRgSK5BLlGmDvZg45YHS/vz2YxhnZvPcbgcfQiZXcMNiQnUYpAJBjIpIASqv
eSwAeZoYMxkcAhA4JiTMBNvsAGx4WZCH2e2ptzksak2QoxiNLytAoUVlt+lr3fqrnFOmijzqpGqP
b97YEr+9yTbYQfLDPvfC3FejFbb6FUM4yIsCBkUnpO7kX9LFqDIgVMpKLGxo+GPiBVQ//BkREq4f
LwARZPMjNsXJUGYyX+w0eUS9c8bK5AHSmXc+IcOuC0s3lT6t4QFqga4iS3UIrvX9vTmEVgZYJiV9
HjOm7dF/rk2HaURgb/Eok287p2Y2a/Ld+qCQaWL/0Z3AX2CCmg7YbH5h2E9n/wnvMiydA6xNoYOt
GOKP6X/9WReuIXtOd6hFemTlhmgjderZYAMkxEB120OWieS9cDmi2+u51rBQah5WxcqX9cdD/KYv
k6D1/YJO/ByPy0IGvehPTzl0ImMRZbs5ec5lagYh3yVHYqNRwz0y/MoO26ZeKJzlN8CLtnw8kROL
G1eo9PuuwT8FAL8ziCyjF2JhVf5t1Yygb8olxvq37yjuWRfIWWFjYxdXZVimVjEJ11kqcL+aYHYy
NPKNbmVgqJR9H4v1twHRscfriwNubA3bilZuq36qq/8b/ihF6SjYARuv9TjXCuvxu60i9Edo8MHq
NvnIrfklSQe5dxjqECOi0NIQxkkbL1at9uhszkYBxBuhfmlxymByb1PBG4Lr9pmUwqVJP+ueny+j
WUk+E8YOWyxOm0wqUGgtfDXxPGCjso224YJNfrdSNL1GOrkqWROREk9pbbefM/7O92d40QHC2bLe
9Gut0iWP3XZRfVv+GgVFhlGE1NBm72qscgiqFfWLUd/yAGq39kEpI5oj9p9rzw2u1MGmqlMwxMzC
dJlh2REdqj6WY8Te8PsSiE7/sFhc2q2XnNPqvQF1b+ZDRFe3DrvenNuEOuHsT3EuhKIYd4UVlGAk
Oa5EjqpCCHorlBV/jLR9e9qJ6vcenjU6OnOzTCivm+zPRmXtvRE3rcV37Oc5B69jTwavf+fVo+VK
1regnTsSrVK6j4ZUk9ZKEFYUYZgd4PdlsNmxQBMB8pLD5TsNirlBXhHE1zzs+iygi2tFxO/WkjX/
XCGdUukrita/mmAU9EXyvXylMQnDnQQBM5Aa3HJ0D3/vw58psaVbq7ugEvufkknBsoUYlK0mSxvF
iX4fYiFfxAGSF5iecgfzUO/T7R+XxO5G56lbHAat8Xjfnaz7XEjPRTfCBIStYv3Wch51YPL7ce7V
XP/BAUl/Yl8bEZG8AemkhSKEj4tXCq/PYrrvZYedQlFt+RW9CSPZA7bwh1dk8WO5iBQnlj/vJph9
E6QzgghoS4oAGcc7uWgtTcC7o1IwDYPuNLirAF+uumFhLJv1B2k8/QkX3cG9iHGyAUwpUrDj+ger
ZeTmcNQDog4eT7u8LcJUwdUenTz3u4Dkccn5ry69hc3LTk3x01Bo9ciflICG57OqOIEimKE/0Krs
/5dxmUmuIzUj7digVIofbH/SsGjkVdv7L1a04jEnRS4UJ3FqOS8aCihQ60kVN5rEQLEMbLsIeTip
VS7qMpYBuj14qr0nN0jxBC4ONmaLixp4vqNm0xnZ5X0HmygLq9W3ZXVMOvHhAql5jA3tlbDnGsvs
1Ehqpr4jEmMHJivgb5NuKL5D/4xRx9H7JCtp/hUfS2jKfDJ76UiiaFoy4u2fTdft/eN9J3N5r+MS
nTY1mnw2yP6WAwdyUMiuSsCpJ+hhMXtBKqxYbob40+R0p+7oyfJON/9TMEDlBidKhHXoDwzYJ8no
jD5UXeKSCBxXrYO7/+hOBrHZ+i7pP+8BjlaDlRSjSdUUCLDRL93Mnv2iawehJXOOw9M5UJoHfxh4
ZS82xWSJsIsCflLcjmeronVKkhJqBPYO4nZFUSzcLr0DfuGGu24ZwdtDk1WdonxJPnsup0ho0kOy
hoInW7MsZvU2oMwZB1ktRGr9fXHoP7YjYoWlcl+rXzcruwV2HCaZMsvIYi8VSRh6T0ePNXmi2iNE
h7t81+U289UGsUXz0eqrMQhzD6jE+N9WiXOutrGDP1E49uw/E1MFXOI7c/CaQI2W+N4vhqGfs2xm
FlGnBwPE/WqV/ulbSQ8HrP9ktm0CTo3qroXzliRG2Hys1OvvG6xyBQVdG/DPuTumCgh1PDfhO5i4
57eDmUkhmR9EczPA9yI9m8cLuNFK9jK+/S+Ge2R325whWYU0prwq5cAOkShhB8Cixh9imwjvfMJA
650exfH9DNFf7tuh1V3TQ4qeBYn5D9CHdplOJjR8xMdQUo3LnOFcfci9RT6TtYqVtZQOjZx9Luv+
DksyK8gvWUzXc5DMlxUSpoP6iQP5WWLcFjHOBBUD6izaLATf3OKkL8DGDmqdKIzo5aOYqXwA8Yse
6YioxjolSOKMMdpWlugXgyQ2zhARMK7V6qvjV1pqvqS7Mp0Ug3GCV3uie6iyP2DB6loaqp8ricgN
Jh0LI3ybgs4m6SHqJEFxQYUWs8ELKmZiLYgH3BTlPDNkW5/htR8a7liq887aCA5rJKsj07bs/gGF
f4oSJGFe93zo/+gBl0Mq0moxzfcn2nPrr8Q8BMJJUFqgIcb105s5pt/MuSnMikOoBjSxpvZ7rZve
b+3T3Nfssp1v19hmk0yLYj3zeQEPl7+wNiWg//2x6un5bxZ3x6dfqi8X8nXe+88xadShs1H5BQZ7
P+d+gXbP8365OjbmDlctAqVFPfY/xJ7OLeDGS7ddLToBrgz6C0MgncmEGRRSHcmQagc8+4WtI6LA
p8Bj3BaNi63MWlOY81sFad85OlzsNNv2iyGv/mM/Ils6zKn2FHnmNpLDzLd4z7jXqOmhoQn/UZ8X
PZlYTfG02lj0gFQfnLdwkZKht/UNLjX6Fbuv/t2SyGZW3iXhiGZ8tUN7V2MZ+ub5OYD2WFOj6oo+
iqLm0auk37ZmbGijG5EDaGClkha793L5kQmhVepMEPv0Wd3hDtH65qQKIw6eTYZYfF7YZwC84n32
KniV5IrTwhX7f9EBUzzWUXPfkohbjZvnRXwfs/gwPYVzUABmJDfzfgwjLWDvcY/u1pSk1kaoekY5
g20+p/AhwC+mu9jfYCHRWsi775nq6Kj4XtntrlKaj2ah6rOMXD4HKJHWSXwPYAtf90G2xyV6ge6m
mnnabpiRhdZMkpqKP3oKJa6bsr0T3vflG5AyJt3kTSY05VOqXm58J0LKyZeVtOKqKaJ4FJoqC3JZ
wsavrQYY65l0YuIW0CVnEuigr3RAMSFfQC3oTaxoYauclHB8acOeJgeBniDtJiJtakGISRk5EG70
vCgvj9/Pfy7c4ImoKAW9Pth4DEZNAkXQh0Y8w6cigdx89KX6DqIPFZmHAiurI8Z6uvE5Sv0juoy0
UetYdGyxnhldzWhOwaQcod3AdnASFRDoliYCdMF5TOEuJx/fkrvX3UUZyQ7OPdLGyymujn0PQq2f
t4kLdclOudpin5TYkYOpH8ab7P9PDXjEVoc4s3PIzJHVIw+qlb+K19lOAczfUDh46IOkea94sDAH
2RZMOxc2FG9KZwc72PpmvDNh9+yx2/sRi25i59ePVTnWhBUWOSFNJmWBhvZJN/TsnUKe826F4IRR
v18NFFvw6BEJC3AhlJKLqzx+L1R8RYLxqH1oUucbpbhupKO2uRZy3Br1unwf+Yh88osxdWiozGZO
5sVxjDZuPywnHXUKl0v+182zvEgRXl4yE7ivBL1jUDy9MY2KGyeBnKkH6Lhf2/8v3e68p6GhZe5U
qKt6KRq8UoCVai/RNil/zRAkcuswf7jYu9+uo8rmglxBXrY2IP1M+m9pAh9nMAgGcc+tCXibL+eH
zRpolTu4qDg4UmUuTyzpOIgWPhiPicISyq3NhKyEFvxAOrFdvGD6+tmf+WC+bXT/axhUGpMxjYey
OEwjxrZwHFKjddUJ2zcVUuewjP0I2kMnAd44vPFB+kjE9SJW2lIp5qNSndn6sVgg69ckDQTAWhUl
dx+SUj9csyX87Z8xXLHk3Sm1PH6gIykTISpHP8xC7vZ6lFBTEaDvIyQZ/hGVYYKd3cd19dAuuBMV
Cy6DC/RpFMwRUcaG0N6/0nMjfcpJAtqkXlve8L8jsCR00Eky3XDGEygvtJ+TV4h7+Rz0B5rbshPg
gWnaI6L08ViNuyvqW94oefzmctOuRGwNBA8azzyWrrs7XMdSy6w08B+uyWeMtctY9jJjV6pD4FHI
bQMpvCmeZjarJ3yRiHg5Llso1pmU3V3sr57cF27WLdoLTjj9DZ/a/brZhDHHxvISsIhw74E7Ux4e
T8LWMSm9fgfnx64cjvUqqxjtAV+WH8xIQWuHXvwv/SZbwi5RkcG6DhUg93ewHGkocyz8iYni0m2N
aY5O+B1oPVjvV3gMJ5uGeZ8DVocoTTUYE5U1YUygkvEE1e8/h52QzQ1lbjO05/GZnkC3DKRWcZw1
59tkmlxs9xQZoEax4vbPEBunWMAB7yLQ9PaO+MaJue8Ta2DcfprEONaGJ9EvBLknxo6w1XPQ4wNy
f/dpT1BDTlhkRc4H+JwW48FqCikW6K2+gqQgJP0He4wnpK+kMItJCqCq7TeV0bJe83a8u6/jahM2
60L5ELitIglOIBJ415J0XDq2NFYzGuon6gqdxEmv00XP4i8uzc/MIqCztomzRi3XhKa/wsKT1y++
/j7A+0upoYLSoGYejOlIRElokQvI1t/oVY7ZSLjd5rfb5c9xHeRY3HetdYZCJER1L7623+28SLn+
xzbhFCEOKGldzR7vhdBni7Wdx/OBVtwl5jhoOnvplvd9aJsvWArUG0vwN9kJVW2h/mlUEKYEF4p8
pDChVM8obYLnxz67igJZv6HTYavNsIpVjnHdQ8Q5jkV5F6pbEXM9Zyoe5gYVgY4SSeAOqeEKu/vv
a6E9GX12WIfw1DbLyUXWPHu6mf2bDIaefhr/cwsEf6u05Bne6sHEDvFmsZC/R4U3qh5dBmB8mKT9
laWnHsy/9SI25VuOc8oG/AICCW68XKfSytqxppCXFKDvLzAImaOu6c26F50gWEImJWrX3dRDyM7N
cYWmGaZXO3cV/s8JCJ6ZqVXW3tVrzNyohSK1iXMy6VfHtZFJQjQCedP8MlYlPLyj5zku6TjlB+8o
/yNLh6XXTsBqpYV5+VLtmZgZyLgCI1z7F1XwOSrLeaUmLuA0DKq+9dm4RY0J1KeZkeZw6cNqKgqe
by6aSNTbNHG6VmiZ1z0q7MkunQAx+MLl1jpFlIZf/4cRoIaRJK+B1aAzfPBzjQmgD3+zNUm/fPlX
wq1f3MyHxz2olltvOG1ijT/qETv3wivT2DgWrLeJPxJv6CffWNvcq7NssSo48pCvu+LVRvU6otV6
kZs2ytD5TNP2x2rQG+NkhkCzCSJF38mvFXZec3a2ixrBQLNpjYicb9Sl4qN71zijKXPwqY3tP04m
ldhj/rzKdO9SRsTQr+P2GxFRuwV9ZHkcIKli98kg9SCXgzEs9E76LUgjTDq7v4ISgkuR8Zles/7J
R5zbuWyUbBca3yoEKPJ80GU968OQMYWmGbHTbdiBjAmGbeL+HT18PFvLdZ5P+KMwWYbOeoslRhoa
Uz+xBczLodexG8myqipI0LOfd28yJcTicDuTTroqHpNG3KFa7bkWinP9HxFIFbqvaE6EP3ooTi6Y
YQLuhtw8ikduijPBLit0Mcnqp+gUny0qSV73VXpXvzttSEJA0w9w/dmcUE3oezdM1DwerPVa9TRJ
nTe2C5hom7Gr8BYOh8d/dFwgUOih9qzT4KGe2IV7Dvobhc3KmiqStVkWPMUFTWD7mTtGuiRZA6mY
1gU3fDsc+ODSW2hG/ooEyY8l3Nukom+QegNJUnxJ+YqBGIdmuP4ksK6uXKwTwih+0ZDimqfB3ri4
wtp7XV6kx+4dW9uJVfHa2mEPnwjUbDK81DdvZhoUdMesZULm0ljXl+xMYgESS6FsDii6FYQ5Qwlc
zbV3j77pH3R/7Mhc6zaWPFirKrYWI8kpZoNdIQd7Il+kPZfU477S+EydZ92U7/sXhr+yPm6tQsF/
b74UbxMjVx8fX3c+pkVF272Nv81WpcznJC5ckwgDyuoTB/5vP3lg0dQThEgbgJmBB7D5KPhOibU9
s71hM5awX0yRSdVR7+8VSgEYyWsfCn93Wd4xbjva67e0B6xfPMrZSzRnlGMInDDcoSZ7lUHKeQKR
3SGtRy81iBWrPB/aEVGj3Y/vvoeLNg3+Oepbc+UZmgIzRdA/FpB1uF34gewjEFNWKNkyNEwC3ASb
YzGWs4eJbanrPvFcfmf3MpbjsAjSCpU8pEhlJerI37XScRbupOQ6/eGGf5VCRsvXlkrd7DrBUKiF
LQSxWYLfkt1bJMMO/cLfbhGXh3Ses6s0wDf5Zvbv8rSJgJvx5PAjhf5hYLbCkzNAGOW2Cmqj5YYS
azEOhJZx9h0WMR5/e2E5Hyduvc3zMyjXXJ5TcM659YCuWZEvf48Uf0QtQ+lEL/YJwSl9MO99UV3x
HZOw4SzR1wndWP7tHQTunQK7DnJwUemnatwQIogM7mxqrDVci0614tsWWVZvhtp2HpYmJ9z20b1N
ohuJHJlzT9kedkRgBlqeUVNz9BpQWaUGL7VKfVBQL9ohsSbZGsd/bdt2eouBS6n8w3aTxl3bzcil
XSWlNkKudfAeWVhIwKl0kmTtEciWzxiNdKHWb9btvcAKwMQmp9gw9bTTfcPxepLLpUUBsJn55v/1
vG3LgNSpPUuofwbDTBxT2xoB9Nu4PEe1wx+t/CiL8qcjoK8ARfDQUgbs9HxS20+TdYZklo6e3RlN
2W1XPY4qcEj4ZsqYJuZk0VIPdsIdztaHGckO3skPgjtr42QEkyA4NXq79KnjdB7ntCNOQ+xeYDd5
UdsGFQSyBDvv3Xx1nf8HbX4wKhce/uBPb5iHVL7N694VIp6n/h5JVv9Qd+cmml6Hl1H/zYl9XyV2
y1i+LP72jZAq4J2r03AeT51HMCSnFs8v4N8cRMlUQe7C0u84UYRTJghdJZInUNt7bi0LieZDF2Wl
mne4QhalZN4THv40iuaIRBEyd8X+VN0TV/WQnRG89RIj7UtQXDhbwXCBZ8R4vyn9jrarobztKbTJ
V5nugOGinBomi8GgTkFivK4HIFKp/9PRcyPnEeaH7DKgcH6Q+dtc6m5WzBMjXh9YTd3AArKcdDYD
Eg6nRvknwvHIwEOgyAjjqft/e4DZ1Q45lMNBelj/fzCgGgWvAX8JYniTjsn2L5NSt4rQNS90cuuo
xDzWfi34eEM0zTk7p7L1SO2cDpBXPMDKVqgTRnlwbN7zqi3byXN94fTonB7e2gJciFga4yQRvsY4
I8zLjnQbZL4LbrUYOCg3dSNIaf/kd8j0JHWmmzI5R/S8IC2wtsnxVIZteE9PaJEguHUjtYxb5QIX
TpIQWEno8/arbr/SNho6bU8mi+tyCg9SMBBePPqAxmG5abVrl1n9Dc94E4dx2Mq9aqP84kvQakCS
mn8A1K1SE74sZcHluWHVtTfPjOz5q2uIEkg9kEOSsSSbos3GJyTJ/ebNDbGS2Wm4ROk3Rti441h2
MXVw8Mm7GltDjTyaaaRklMxU0Vbwt3p81RXinBzRce1KppNGRIuglggekiBRMYO1ACa+yShFrbrf
0AKaXRays2wy779QAlL1xCGtc9Kw3eo7JUJxMFlMqfYuxdAjLxzvKcWY/dJ0LAT6ifkTqdltMv3s
agiKo9VpcCv742lhakhycFoIfhfn6m2bdzV3ky2wYEG5uPF/cFyV2fUZxJgLtd8NH2gyNfRSkouk
N2xdXei9QIVtEOLeWtzo4+DfqU0t2uSye6yKg3puwkAbX6j0xFHj8DPCv5KTiehHKnh0f3FQIqjX
klWeFebvgPkHTdDur8F49BgjNNpLgsOcdsyphpv73aGDfNhMet4h8yc8xDznLDp8dJBk4UkEfF6s
a8ujpPw0488oahFuRquTOZAyWBqcaukdzT8AU3Q6iMi8NBouwz3SyY2WcqGwkncT92QshMH92fJO
70MO0Qqx/6zZNxUUZMMgza7CEH/UwaIATDBJnuSdzWUu8w3uaeI6Lj2i5EzQ3FmPYx5J7T4t15/W
boqjlk5YefgkPlfQVcvf8if0byL5QcrMODPLxAiLv2iOjEHtvkDucL1J7oMiW3JgqQLpcMtUJI4v
5IKje27rbPU40UWZf6FX0hx7QFBRnBgondc55DZgWdpteJpbKtxb7RKkm2R81+C4ayIy7WI7v+Vh
rMXVoy8MeMfZJqBbIrh2U0z7hK6S9J7NgvawqIrdvaa1865o/lvXWFfL/99BdvqwSyy6LvgNEOGV
Gfx2YaFGBEZVozrNv2FVG7KJms5mq+iygVaOXh3O9zbXn81knyxIEGXILj8eICUhpg+Uk3pEGHb5
27fWV4w0MJJxrK4Im9C3+1v2cDcJvESSS3FI+zsdpH//99Ixe3j8Miw85Zff028Y08syZNyUivk+
mEjMQshREeOI5aX8iEkP6/Omx631KW3i5u+Pf/VGHD5s2T0YrVQaW9CehR3hMliyuawczYazsZT+
5xqFElhym72b6zBFF+Vdp/WJ+Q7paG1pb4RzYIiyE599CRERktTsa09M0MAtBarFAmyW9ynHjzxF
C/WGdbyOugfLhcJ7vlpUQ3KQNIUBAX/NMywkQTftrMNwNQgq0nEKShGQzHki25bH/2xCFCH1FkD7
smQWnL5w0ywaDWNvjszufZtLhEnYWmgaNwddR5qeFel7L1GzjulIcGbO9+iK6LGmkr7ufuT1bI20
hZsZP0treiQPyF0zVy6or3cujc57G30B0Q0KUItSmDQTjf7W4Vl+R3D8EW2mLqXX3iEbuKQCSSsD
RpHaWhRJPt+BEzlA3cE9gn2MqDu99mrWp6oLXblv5bni3HGwAWAJ+L2UvJu93ZK9y5WpyN9xxNoz
OWBYT/lZAMi4pkpturoSekDu5zbgJR/gFgX3WiTzQJh8R9SGvOGu/YEIhoFHJkwZO9VMFjQ/QsKD
qiq1NmWNmf4qqaaEVfNi9uJCX9DV2VQd53ZHaExD+GTQSPlnwMS/Fs8Da2NZcN+C8c9WaxT6lfGO
23eH4mrJInwHSZWA6S8f1kR6AfMsb3kSKAVOms9ZVUYmKWHKUYDQ6s6SABAgwXPrwDLVomV0xOxy
bhYJIfCv8bG4ZWu8XkdZkr5tFeRfaGwLUl4y3K3Bh/8WiA8QKgOTDpk0ueyC32ErSS06ad9l6sE0
tX20L5kXF4tAmx60NE8sjmBNMM6s5f4iOY2OoU+XyvRGrAPnRPWnnQg6nlPGJVdAqYtrOSs7WDxy
xJNqCvPavbTQrw2ozdynuE2iDsx/dXgTP1fcYNm2FXlLCA0VgiuDXR/VjH3h7yGex2WV2I3oMjrF
ZJoeYduEWnZ+37tB/cXKm745wlXWpW1HZB63G14LdtKcV9PXYJDBI7DwN3OOL9vdu3N1R4qPPUcS
6LXBOypDfhepMhpBQLAQq6a4Cfr19lVtKFPeL0mCs7G0sWN1Mn9kJQxyI5FqpwwCECH4PyMlcol+
qJxwvETj8Rqnvsdw48vNwT/Jt2AeJ8I6H5fHmp5U2lrPEmKJIoQEd8j9/0d2a8KUyIHS8bOK2VIW
ycjpHiqvaVIABGXs3kRh+B8eS6TL3bGe17MS3Z4QbfitcmjS94tExxtG0PlET2pQwCOrnsDYQWzF
H6x68+lBywPro5sNHPDvvOmqbkf6pz3OqANKXOZr8S5i9PInNioPkz2DpGScpreFS5pQNzhRZveA
70o/Z1iIEvZN9lT1DxwxaJWLZ36x/1m+B58P3nSc8F07EJKKvj6rGBfnZIkW+p22NqnBv3DCnY+u
/8g9NmjgyIC6rrYukIs+SdfGJ6LBNEAYLU4ykGVCp2AYiNuAi2KQoJyvvM0FCb7QG2eh136hQAYM
p2gSFTEI69XaiapHeQI9Comtk1Dk4SmBvy2bZOgWR4Y86+JdGR+7UfKcdkhThTqRjebSMos+zA5U
Ki74OcaKspkLQpR87BUDeZd0JjOIUGyNDzf0IZp1BJrT9KAvquWXqncjt2OOc0MMCS3/go6akbIM
7322flUVTRChTIn9AIRDvGNy7p9LwafTPLFX1x2ymBbrjeNWac8cytIR3tTR6GkziyrL4dnzpuiH
sB12eLr9YS+Rvv3Et9D8DPDaZshukgOVJ5WacgElm+G5v/tQb//IaZzJw4EFm39FKn4u1KNKVOR/
15rYpOVimr6eoQiRgqpB30GVr1Jlr3i+SBGiVZUchT9daLdEF3JAxz4NkRzzcExXyzUfOiZ88uYZ
H4h6Ca7x1z13BePbKaSjZsgIBC4u2Q/qtg1k/ARS+r/ZLPGrqX4iA3xV/tpzll9ojH3fDQcIM+jH
jBXA3eoAbWh1ZD40AhVIGONMO8X6hmv8rRfhZ7uoQgSQVRGBJtRF9Hgk2wHLaWRjqIPIkFiSfE6c
BXcTZss1tDMBrqLjz7YB5FhNpL2D6QxxDUWzvalsBjnNbGHc7IZQbBzUIEQyFvxK4botlyeaydi5
WFK6/9Fw26Z0eYvYLZsDr8bwnxAhoVKcSWye10+JULjGLDSRP43THZDuKhL0wsOKMNAqjGJQG8iJ
67AoI4CM3qoH06Qs/ciLCrmAdpfxcKAUHDpcZE8Y+jvJE+SkeKyHJIK5xr1O1WB03OQ/hQ5ZI2Wq
LgLmqBo8/Bgbs9yto1iiSRtQ741YprOTwvI4PFAiVLT0u3xwifqf4aQOnOkaF7dr/9gYf7ikmbr7
UAPOQ7HAU5rLestalUrfu5ho2Cmo6Mu0nvSNqen5Fyo1XnOSMVUIw6ZunuzuRgh7+d43jJSpc8qp
/ZUTfVTuMlg0cKV15hVhrvNRmqRJd/c4GDSvtJd3k/QjboHROxePmCFIwrMeqRjgg4Z2nvpnk9k0
0Zd8PNo/I1you3ZciULjsfpLfG/DtVXCfmW4emRog0naaDnp2KU/rz4HjVfBCJgtQUHQAzac0Zri
za2TcXiglVhJlU4adjxx2J4x+tyfS4Y/t2EW2kIGl1VrEo90JE7nRewSAIQkPggVpwGslsfWHe/p
bK2Im3sdO9bEmjqFos2AgN6OrV2RYUU5sNOpbBeJfRlXRdZKsYYyyf6mrlFQ9QgVL19VzDEX+zx2
v5OegH/pA6O6/yMo7KTTPHvmyasIzT03Mkz8c3fW087180kKtDnlhD/2Y7BDEFekL0DobZRfer9o
SmkKdli5IfnVLrZWbem+TrzKvcyg8YyL8N2fgAmNpLGUV9ibwFBcHKuV1DAk+6Rnj84b5D0A0ObS
us9rr43pPVepBIoxvVi6HM5TR8DwWoir+PLRUKTmUj8Kv0ANNN6tz/E78cIc+iZUcpirgfnhnpwL
mtOS+I97YZ0S5GkcmcWYl5MYf4De+4KG/N51rel4V2sF6vyBSV7pYSJZukohtui+FYkPmM0I23hk
zQqNLd7a1f5EeeemJU0vmcpBP+phHC5+tyCI6VyUmjsYWFzCK9i2z2gIij0XlYCIWTtwV9ON5pc6
cdB4R355AS0q23JLQA5UutAmTTKqhdHSV8MtQ3Lln887DLD9hPM/G2HY7IbYx4o/1StnET8FpOT9
SpUbidLqJvfWX/AbASElr39bhiHmA6HXCIW8i+sbCGHpz7gKokz75Z6IAyX5MSOYSqczfdEspDXt
TIlAhx1wzBTAtekUxbRe6ZX6eg94L0eOKL8yAmeJ843mTusD/Ab3HG/FPfxlUqFR1Osz1NG/uwzi
59QPdNyTW5gBnFKNqpiELN619AABl9ayDAelYEYrDPUDHxa+Gkh6KGJbLxBC4ErwUd0L6iFBnSi/
A/pi18MY0e0lSX00eVU9KSo+Aa5XJwKBg2W/8/ifZUzXOGKB414FDl83/Phkj3wOtZvSzZBFbXkD
9iyTsy8D+SXbO5SDtMz1O4qMuRlPp14i+UkvI3AvNmxfDrV62RCwSHDlyyPoJsoKMJe2mHnAS4SQ
IxWvbRaBWSNjGr3g3iGXSu1EQAnIwyawSGfuK2HZe9CtItzJ379zjb5AGAmoSqPsisxtwHB3fBrK
/vlEdHjq4k6idXlaBkZUulMvTwwO25wJk2bZgEiBY/6kjpXo+xabek12KWRGz0NMBKp+9nO1stxR
gRAy+8WFUckbbfPlR9emVMgPiMDazWmRl6R4TyMDSVj9nQrFO9ij3oiULYj+JYxiig9Exk3Bn63z
HS4JuWdQNdVzScAHBaeuwj1+BsgdRbaI5sBmfZu50ehKBRuo4YrMhwdiiNQNxLoreNiHfxpq77MJ
uFsW2qe8mJ6MVFFIiGQY7cdXmgx4eDgHIDs9NIZ7kGZIFw9L/Iamgge/SDIW4sbm9yNYiezkbYJN
bS4VtO/9j7fMuprvzyVhRjTAiFYcZFh9tfhgqieyKYSv0MLDCzn6Isx7h9sP7JTvKy7vsPbWXQ/H
ZtQDLt4RBSNuIDgssirxBtbTsxpZTZn39mTvxzP3K2jOh9EA3V8RZRit+ERofpfS313oemvb3X/Z
RsBoc6IYXAkMRSnM/Uqp6Ejt6CyLqrvCvWR6s3NgDChZEu4p+ydLkkeWtH4jWMIrzRPD/lo1sfKe
1xX/raqADiMS2i/wzo8wqJgKl9gqjNWvXF4mgF/MLyIUWbMlawDx3h/IpYURoyrms/Qju5UL25x2
E621qqJw7rPSl4MjuNOS29yJdjGpbPNlAMg98M+sgsYkkhwaK3bnygvcFUXCj0ub/9+guT2pmkBk
+4knP8U5X0MRIW4y9lTBq6InKqJ3HuyH1iZoOdgFtCKJ7gwkIynitvRQQP0NzqtayO1/D8iShfLr
aMfpUkmu/DO321GLhaRbSydklD3Wo2KLSWRoHs2bQ0KgCT7UgA6N2H3SmYNuPgRTXY2H00gxXoAy
Iv3XgcaWBBonbJ+H/73GMjlFtIadksAjXNFrjl3cOlwYKOkOR2y4c5DUJpEboEPDyGI3WDrVsu1x
DHGabYfLlSRtJNyiuuv4yYHUc7X0voiRIvHbykQQAKrZjj3thmYunHexucvFUMCK9AkLo+22tzeq
GAn4Y30vD/Mb4M0I/kYvTl4Ze/oaY1RQpOPjq+XlAWEgMOxhitqb7MSQfCrp0Mx9gY39Xh5WxKVj
I5DT1Q/XdLVMZdQQ6IGNBlK9DFY7HQXpK3zm9KU3gRhwnE+3Y4ocEOSPrvmBZD5cAIb50jGn0KX+
ugEiqzm8nOEutYwjY2VTXqf8dbf0PVzRLRv37OjanADgFsMQpxq4aVGvUE3krz1DHeAGM1EtqRQN
zMx+vQB09ZozjU8zEzImDXwGes+UHc+/1Lpp5MKDa6KyQG9tmkoS55TQmBHai+Xno7JyCWBwJuH7
7JC4Z2PvDR23cr2OAMYv5ieNUgrFed3pMnuojSWcDR7hqFjcHY4IcGEQZR1quf6+UP1ib425lPJ8
eCVLpEbG4C+QuxucN59u+jqg79BEAPydq442TU0eBAU8zDyjK50cUlaC9HXPbV0z9PgCDLQKYzUo
wLjsRkH/6xdPFHz83Wcgfn+sxVgrDgdp/Xw0yqZfyxAgCTx3BTxy8s6S09YG48ZYIVcpvGubfTcB
RDAgpd6IBcsaxlAhcBmxiZN9urA0mpuFsQOj2BnqvfklQVxG8vzrVsGg4LxA9bvuyAwCS0Ndcu6x
SlznwKCLlncIZarVv+oOAczmQHWDMAgg9R/Yb7vim2Imyjfm1T/tNeIZxFyTCaD6n4WPQ1Vkb6Iz
qbQUyn25212g26XZF0nFVZqo6z+kr4eZNZaxUfvR1sae9mUITECyuDFf9HGoToFcv0vCV7N1nYpp
TGKWcFSzylMGdiX9gCuWmgsPlsdERQ4ocTqwQb8RCBae/y2lYwrieAcHU8chfa0Wzgc1DxXBS7vF
34m+AdPZ3rYxyKOzNKefFIiHHKqenEuDC//b1sj0cMuewnzSf6Fz7dBNqCo/B8aPnXQ/x5Ry5tO9
ZnlOrsm3+rm+JO3dXkZ1uE3ZKowcjXIMGeV017iteinYQpSD1yIM6wJxM50jRvHn5ZkAN4ciTvi9
aGeSu2bfxbHEMt6RGWfBfHx9vgfLPbOaEfy85OKPdIGMHwENMOKHbMELFiHcKqmnDiE1hhtyo/hc
OJijksHgldaYtBq78YLGhKxMFJO2qzauPUrSvA51fmJ5APOUH9O75c9nViweuCnWFB0139gunHt/
Ld7TsI49+Jah/kXjBy49ouBmqLaCOYDuGTH0Dqzs9TS2JR/jJxE+R0SP0hNaPWb/UuPva5MljkzY
0+SlhtC4eEDSY+iO0n3F5sYxIyuzoVO7n0w6H7+9+F9Zxvlxn66CX0F/M6PXb48By/aiTbXulX4/
IpEyKFkK2ZzxoPXfLEc5LQQhVfpUp3WyXzqHlFQBJXhVEXLYRVxbgsBWK0RD+MK+d1LjnbisyrXV
GXOcoHwBi6Hx9MNepH5mwXguHd9Z+O4Q3zaqEV+iqoa5YMWGZaHt8spl1hDMGxsJz/Boelsx1UwJ
m0VmLCU5Q8gt1qYg3LnIQnW48uTkz9kA7AxqWUF34pTSMouaDn7+ah3+xVkERSnzjtfUyXZP7c4W
rytWkoxKwn9vKk0100OtVJ8zTCQUSNbCGjKL6L4AUBzt/pXXUvAUnKm9R1XyTqa8SSPIzgXdMesc
o5f9+ujQpuqeI5DLJlOtURFhknwNLCy+gNkrEtbG9ACuwgLG0YJAid0v+bdJmCfxrdoFVJrnp3ZU
57Vk6L+VHUlt80V3v9q1KKC5vvYzq4Yj+LuBObmcqo2XtQYH9iMHBVovhlK2cdWvq79jMctdWarV
18OnM+OQCgr37jePF4BawRACSxaZ6BNQguvLohJNGLwZfjuC5sUNI2dWewVWZJFOUZALE5XEKqKG
m3J3TA0JtpKe39NhhpnWrl/VfwvuoaKjufrUqjLLwqMGGW8jnHMH1GiwWdTwP3ogGe3axaL99KZX
yg4oXYYt4UvwXROeXheWVTd4CdrTmFidmtWavE9lxdFa33WGfzJD4aFa/P5UbixJLsixMO+W9ThL
+gso26gob/meuCSjr4VIfPg3HgOVUXH8rbZ2/NXolIzTaJ3WoA/kpd78UortDNDg7zJHiFjDBA7Z
1Kezqqj8W5EyxbtV4hdJ58C/onx/ELWNown/yh8a23yPrTNAU2BJrDsEQvfwGkBZgSRBBrVUMTVb
6dyTZ12RoajjiONeZy5zAfNU1EJjwnfKdxZI8X8y+oVDgaNqeOnCPf41MwuFKOtvUZLuaRp0Ndxc
Np5kwvX3as0/HZDAKbBT4Jr8spnrNU3dHcUZ/oT9A0eKo3NmFazYo4RxKQQlDL4CI70Ts1NbRBt8
UXREur90nBU9YI7OJzQXxUTMkDBCmue/YXdQ0IW3+XWAjIFvwwSzohMAflWeM8tCaVRiqYW9bIJ1
uvFNVyVGT8r+JzMqjhcj2feOXufIilvqHf1MonJkhBbp6i2om3t+e60Uc+Vjy6a982aDCz3IK+Mt
c/kUT2syZzrf7wbZSO84I1h2dtwOlGM7e6ncAHVEZY/QvQ6CVmc/RjsJWL8uDU3Xjqblp9YbzmP3
Sm4j3pvd8T7aXjXrovIel6TVf6U3eAw5zFhTk/e9J90PtILfJzIhxTQvQQt9D87nRLxCNct4hlR/
iu8TmBdXB5mSfblsiIeFolsAca5TKoaTszTQEKlTUcq6oLF66/xKWQfyRUjhbeAfTKQV9ZqSU2Wx
6fa14Pj9nSReXecCZUyQQyjECDoD76LIlgNQ9E9Fi1/9Vli+L9oSB+FyjnPceJm9RW32VQAYrjM1
SKw9VRpARORsESOYCeH//xvEyETKyI/ZN7c2WdcYZIZcQGkHbsjdyUsRqWApXgIcdiNbTFKRf/Xc
pCxg2swDouS7MMaKzCtV+EsCyWEUElZbG/f8sUiP2xVoEh5RKiSuzV6KsKJ9fEBxTD6pDWgxmDVj
2upsHaAcbw55dPJRKrR29ITPxCfTuaA48X8GsV0qJHIfCKxw48bGZ3x5tu1w1iOynja6Lu+ROznf
ic5FzV+TFFSVbjT8xpVBjfX/JYO+czEdFk4dZvBx8nzCrRzI2ezOpQ1HfMmF5K3mYJNR3TQq/mDM
iwPPiAWdgAgr7lJo2AmehI99t1+YI2rR0idZB+fpXXaMCUva9I4XCZNKk2vEX2W9uhAT5K9lx5sK
DGpyL94jQiZAQNc/VhmM2R4xWl0HoiDvIGE9A2BAf1drkURYzK0rvLr0EUX60QN+KG1W0MSOxyWZ
8MsliY2IAoG1O7QCT/F4HzpTugRKkTbAJNnxutq/nK8bR/FYCymYLg6cayM77nVip9aovJ8ILxHU
zPx2pWKdLEQr9/q9kBIZAWZ63eQ510R3L2hyqbzg4sdQ30U6pvffTVdft6b+fpiI/6ZAF2Nn11B3
vo75+AERw2GA6Q7NyUaz4eAUmFTNnGEn6T+AiYCyp2S4S3XM5bLDumPDwE6ER8eQawfgLYsrr7j2
YJmRRDU2bhcwcHHV8E5zLxyPtbMEzDoC7Bpa6aOHbFtCUXpadeH9TndzvbKWAoJl7IhHPefkCdmj
1G0iJ858Efz1lfVVU91HrHZDWtmAB4bCI24ZGqlhIOEzjGdsDuYjLCJHrERZwVuFfy4mSAhNN9gT
d3U7lCBFAK1x8wBlm6BhaoZmNOx7omJg7UWsN5T8h52g14nqZlsSIYfO+ZJHA/HKIIrRa4r4rP4g
3q/9wDq3f+kAIDUmDxzp9LCbOW0qaugTW0gWTsOmSYBjMpz4fpogb8hhA6OVsGXvs1b3zz8LxxHP
DhbWDELnrT23bblN2SSM2B03Z2u0GlWAV+HTm8b2HiL+xQP1DE/Wfo7X2rfsgR+XZFUQchxDfXTr
bjFk3kwDD43wbsnORN05zk90XfB00b6OIRl1GFdnBOEPx04u92qr7TSbL29L9Ln3QWlw1oS93DVy
jNw1IAg5vKJdpuOjmoCPw3pc1WixpOUjzeXq/c7t0we6lZrIrPhZNcvzVEpb43WAoFkcwHomAIKF
ZsvJe8EnZeR5hPr+ordsdM2oAefpSezU0ne3XEuZ23OvUO1+DoIE9LQBKvLSr+smilCzQ3j9jorR
zdZZTHk5WiVOfAsN1Z/JnpKV6xKMHYRCIBkwdSfxfe96u8ISvBQxTzQFaRiTwZ1/0ZFUqdC8qerq
vUVyx91DdYauS3/DnJ1f7oKdePY2RTje1yka7awY1sgwRyL9lz+YEtXuJ6PKIS23gpYT2Q9OXf9f
AUtJI42Eck7VdjDwkyyGpxjto73adwPL4OwEKXo9o1Mss64d6IhIAucDwXsa9r0oKez7T22drN8J
GEqi1X18juJ6PlENusZmqPbTH2SYH7CiG7q25FYPZrLRKbLWHW6NHkO831ySH0HQ80hfnoocGxWW
inIqMrwgZVtT4/6C5A+M7UOSZjV0f59almU6DQc5JyH1ZqasESjGfWbjaJh2dCpQ7upxvC3gMn86
//VZ4DvnY4cqbWM5eFRx++cuLOXxeh11GL+ovMhPN33sQSJiE7QcIkWU2uyy4lE7YoaFLHqzNbZf
gBwrPmgPliZ/LsuGOFSIgUP24vp0QmBGG2G+HLwjq+GQ+qAylTuB9S+hjslvpR7DtkD8M3YblIhV
k21jfQFoyVGbSvRGv72XmRgXOIGyQvoDGBJDG9x6bmvQ3wit5br4rQmi/NeO9eLWGfZZeyCyEiBm
3tC4jmWOWdBynjJkKT41ddlAkxn1Pc4SPBuoPPsRpgIlkLyHSYFstA4qI73PlCW6V0OLU6/oy+e8
xKCK2PWkdQUa2btKILhPy0qskyjXRWRNQamRNucvBClyByXeIA84tWgPu7YK0JiWpzti/6tOIdeW
GmSmk4th9aAsZ731zlYbikFWBRNnd9WvG2RLjHluogOryDxbiOwGGc4GbfjtJ0XnKVQZU7VMHnvo
LfZWnvV8olLzIoP/gqgsATBbVPrqe1FHJPavIbi8c2PP2O4PGNN7xqbe0nn6z8S1JgzBcDCjMZYl
GkgfY+XqI0/2SbGoAWL+yNm3UcYv9T2jbGqqQhRmmIvxxSWD4tMKUQ0KcLAApwITmDSHi7utG58u
IHpSspc87kWJQmRCHRGmgztNbHnWf2ZuhtJB0iqvgTYjYKDaFbm7DvGMM24w5kAfk9RWRpfK9Dw8
hMFtdpJNlUuXe5vZnRbopSlYeoKTvxsXSa7gu+5bdzz9EEpWz56evWtzGQ3sfDVYT7cK8OWFB9+3
Xh7qPtYm3wlBsqQJaC74t30b7DdD1JVhe1HxbCMiSPixfbLVqEGjV9q+8FiOcycP00hbZQ9fpMUs
h//+bLu0KAaBaAt/ujL8b57CWW2N0XfTpQPv+RhETkIjiS+SdaAGp69Rji7rXe+kdnJKsTQC6/gj
U227dOz0qb2qH3o5wOWzZxfVL88Pt8rlhBpesUrn2cOA7chphHyf+f5Jfgb51jbWpG9vLUZqfqeW
+RXE+LvTOaoO5b3r5KjGTtJTV4aqdx1ySmL7k+lGmiCTTFtowd4xhCTmm8f+qJydhA+Ef12nOINf
Z30FNNRFzlZsX5KQFezrU55PFr3DDxqkdxgHGBpQCAXjt1oCGkWsaFBU5bjHcTMPeeaLxqJirydM
+w5Smu3yPgVfcxbGUf0BneIAPtrk22N60SE2WujOJUpe5F4pfeMDgRvSZs7x4vrPIBBymMDr72ME
N6QzNltPmAhBp+NxNrQYmOcHVHGnzTnkuiTxjel68XcDPUlWpI/EJeiSyFmdVJc05tqsvSY5goZD
j3d+NrMXhj3AyyOPgOeiuZaOWGqSFzfVdXhNMHyeZOJIs6Pb6ZnTggNr6q4jkBTmJhYH0Xvy4peh
iYJLlkMwDOV4Su31EWZjBoDKdQozLaSs8dF5uTnHw+HntmSmL+XCMOrhLRx3MDR66YgZeXljDbCH
pfytCKejhRMmU71beGVfBnJVPjQ+4unlqQR5UVAP7THviMeqFBJa1H2XxQAb56+nU/ml2S8epLy7
Rt4GDoNukyKsblA0UUxd/Wwbj+dVa5Cwj3I4O3G74q0S6DdKhlHvXvwezNM7HejI4Vsa3gOkSGDs
CBF16LktTOMUZgJQkDlD4RV1mPLi1uI124D9S9F6ovyzW9jXmdNGdjM7woxHP1K8xJvveCr5f4sr
c16ZQ57P1AOhfKKxqQRdQOv8EPRmtcPMJGFZ7BlhHLwQ50m1l+BxrVkg2mitoWUPa1FyG99a91hl
cMSZ+RpGBsPYBVQuNUh0qLiUlMtLzTZdbIFHfz/AcfwY0c2oY+FWV5wLh3ZhoqU6M9oVWg0Lv+NK
8oT6XnXH7F4830JgNMEPrVNLwe/Pi0Ylhiif/fL3JfjkttbsjEF/JoK7rXHiniLLloJxaZQxONvP
Eq1HJG6JFnIVL/OoS2ubycydIZQcdWCajFp8gOBU08Gn0GQAP+M8VQfX5jb4CDV8TbbxWBJEpmAS
RU0j89w0EINqSTt0umqxGKwx0M2Gf9q6SWddYqU/7qCXS/Lw8+y43C8YlOBLNCWFp8IB983Maz1/
i0jXcdRsx8d2t6HBNz1zIKeX1mH3P1AkMtkHGYZFLUNQVzscIq4oNOKgx8sm4R69/QzTmBwDYaDz
XCYFw31Pxi6XwERqHVnoQKaTaMqRo8fVU26iJlhxQ9n4v+01oZP6CBOf/pSKPSYhzfWMjAB+YZU4
OSqF+xx9R9k7m7eDqT+rmOQ1Yr/eZkQ2S3F8tkiOqH7pcHzDq7cCt7GV255Dpb8kGqQ8M/UyFx18
ODld26/AdQ8l8BJpTYb1Vv5oTgShnbAtIZnlrZwkGilBRZWJ/BhBgJBdjfc3PmhS0XHxwkNTx1Fn
XRvrsf6i0m0JgCwnZJc7dhYqzfLh+hoGhYqqd2PngAMn+CgprKsCIDxRKCsiQpaa9lYkZpBj1AlP
2h9VIRuZKNCCvB+8OxCKDuTUWNQhiI3bku8l7OLTRMtEFCf78ew9KBV6OjvRtgstRD/2i1Gfd3FA
soLoTOZIa/WYT6Xsh3h51M/zK+IO2gNzYWIMoZiUeOxqPT2dQX1Cp0lsOkqE0c2LUkOQhklMj1K9
2E77a3jXSBXBCPFHa/z7jTV7o8Iig7nK9ZUlf3UzDXM3RKaL/Utx5D26eySt4cDqBwWTHtwe3vuf
YWAIQCYxC6IKZc2/luj7OY+hZIEBTvcTw6Hz+WtocW7zCZW+GWrEGr7RLgEKTyfJ7uNb+Zit8cWa
NYiwMdhKRk7p7qDbDqNLmfdFaSbFxMGkale09Hdu1M40U3VOOoPfPI7lmJLDC5oKr66UIg5gaHkI
VvApHu6reXq3yaUmMLuBUx6yXmOJTR9hd0HMwpnp+aIi3rGggoZCg5OLHXe61XUCiqfJsifPqW+G
iCFn8/c3MC/Hb6H0A3QJXlVvJxF7ItTh1xZ/Px9P55ddxGpmol872V3VBH00XkdojJS+9UFjMqwa
hwKm5jSTEuWwppER1oH5r9YV+C4S67Ok4xgFMu7pqwnuIiDvflDTxnETIIqSlO2lSmKhHgCZy4AH
A+76Klltc0mArd7gsd8cws5TNvLnl7Z79Qfp/K3bkKJicDBe+h6h9a7qhzyZHra5oCWpbqBZGimJ
1Y4Bjweq+3ywMb0W6s6gk4ALIOoPxQJDAXu08nJi9+UjdrYnvygGfvp3Puf+o71z1IBiDDZ7yIPA
a7eVMvdSM6Mxnc6r0Eu+c+JZuhn28pDKQB0H9QtjtOEeAAPSBQDClXbjLTDLq4VMvNKd+FyEMdOZ
9GwBxjpFJdz/Iym2phW3bNLJmex+RReJZPLLYDTuR40RfwGDDyPzX1ox0RIVLKLR6TjN7Hl/JfHJ
+slCOdhT0Y4VzOzvqs52o5QTEWnPlDKOoYREPpkIRduo53dkfED7Y5Qa+TP2xxoPER87vH6DsfjA
CBn5awgDbNwzfM9DRyplwEwUvTZ9Ur6ipDvpqigRZHkCiFEo8daZdds8DzrGzcXsm0ku013sJKeu
UM75Ew0f+5U2F/HUURfJGauo0waBML1DkgMd6kNNOvZgVfU37FAnW5Chz7IYUuQ2VTpIC01qGQIw
+XDHAjcvMUpTqOfTE4dDIp+LMkwsNkDjx7l2B/bmlgqs9nJolBDNU0v8uDN5wRwDIZO5d+JX59fV
PLPw5dXQoQyHgUWZ343xyfRBZYAdGIugp3FDNYd9Tv4KnKoLzEE/GmjX0l+VrBVFzL93eAZV7TLW
movbT6zjsQL5qImkSPoPsHWb3ZWQaRGxMOSJjNu9vHYHgV9FX5cD95mdvgZGgxjudKSmdvFQ3vO7
IroaZ2bE/Fx1FUL7hX172G6S6eh2tjPiA+0KdSVTdJIszJ4PLLlE3FQjbZWZunR2hWr5IaWySU3S
l6OkM8/rrWy+FBTOgar/Hp9UcthAYT3LK+9bHzick1fyd9N2iOjHrKY+Otwk+Dei+hKFiXeIXwjr
dko+PRu89wK8Es3p2WFcv9dzTDMOudSshAe9/Apk4zByCkITaAyM2B7g1sGp5cUrC2sItgHYf51x
tStmtXzjig/VZXZVm8CMaVGvxDoX17HgSKBIyF8IWttsyOBV44sVcidYF0dg6o6UB4EcuBNvSFL9
7W71GcWKOkq+RVb+AO9m+UxvWzX2kwo9vaWwnSbgj5IBxKjxX3vDt4TdURKMSQ7dlSUGcTQ/bBJB
JYAn+DxivEwd/IPzlXfnZYdaROPNib6h4qjOwDrallHIIBP52EUoaPfv5mu7NSEZXeSbE7qg5GVD
vRQATFJqH2lm2RKU+qP4drlvA8a71SYHAuVcs0cOqpNTq8hOJwpXwZt9g7pXZilZ5Ag9LZW27m1W
3Ytppo7j4GQTWdSG/jrBzM693MJORRtLF34VbHDXRF0GavttEMB5prut/SY3LdIRHIS8b9aCzOo7
Kixts73Lx1PA9HRDsJPfIS2SRXqRRASU2ouky/PI7nNOqdqN+5IAkvS2m1+ho0uKrTrANFwtj2t3
NpXCIRZmKGA3iZzX9Wm1EbwaYR9pY5n4owZJz956bXg9XUjaHYWJGL5aUgu8xO4f7yggX0moXWaU
1Uis5acGSItRtxk/kHe56iadV5qMyBOmXI53bQ8de7abaunX6GmoEZh9pFxYN09eFUVZqaKfYQJo
l15K4zL+/g5t64PY3XbW1oMm1RdykJv7b8k3txVLvNJOOOBfHzwkhwIPYYGMGYqdY9yMug2YcAAg
1tLwszxo96C7GL72unGgy6QSAdDGuN05DzAl3bpK5rZBvkLtJ2+1sIaNkZCUXw5da6S0jwQz9Cqg
rM+Li9TEHf/Ovdj6gcteLhl1igKRxlOf5LErL3V2CcO6okT8shDYmPSYCbuwSMwGsW4fZiEYkMib
BMIYWKf1gzq5CYpY21r/r0H2dBFO6zJhJJvaw1VxGPIid+WilQVn2remKasU1NVEZTpJzlkyluJz
10IjvpkEI+07sE8M2CP3S4WaPM+2y44tegGBNhH76trbQUvT3b5g580r2DZ6Z4I4aj/SwZK9tOev
l4JGYl8WZWNgyb1/0fA0H+WqgB4T6Hx8nQcv7BtdpgLPY85f+TYixX5TO3kBies54mV9BBMByH7C
+Hkq2tkLr5EPtRpfMxlHj8eeWhDDhqOpTVxqhdxEaR5HmY3TmsOWDzMyqwWb8Ow2BxHCKVyKMVVg
LkHb4GPJXOmSsO7Wd6uOCVnQ13VnVSGHAGsgI7j5BEy/Ej/0AJAjdyex4NjmI2/VbU6iQUqM89vI
T4Rv00NNvflWhCbuDqdlPXJx9LrY3W99cpL2nuuk32kAYzwTUQa6oYkChW8aZztvCQL5LIfAmtih
v2fZb5YIVhoWIy4Ql7S3jCjteCzWokAaNwDPPRnvtIpoaYwgNAIr8HW7HSzabL7S2DW+oUpV9Prd
z/krasmEoC85a3zXNlisWFstNBxbsrgiE/zkHCIwqor+iC4bf5IEc8/h8hkgKFYRie5pQoQzjb7z
9alfVje8RnOnu6lxM4crswjhCduv6ASEId9k9Mqnv3RH+VVo/x76Jkjy9GWzF2RX8CFj4yXyfh54
t5qBZ05LXVGKD7jq5PJjmkmtw3EnVTSY5EeGVnkmR/iGtrIaG5sQte0vKeIaIrXInvBdYzCR9AH7
FkashYWUZ1MM9xIkbBBMCxa2Uun31yNGMAss+dqVeg2kh7YAeJdjnXnlUbh/IxQuOylWXkBETukn
S4h3hH6+hVCwZXiw/G486jAjxW8JL6S5Sp1rBzm0Xy1KyU21jPh/Njc2UMvtyDgiTsaluEFSprH+
zz2LHdT6v8vJGxm7BQ5V4zzMcz3xxH0dyoSwswTcIy+qbvlZI15k14QtFD8a98DyuOqVYzsH9Moq
Dm+dMH6JH/+EbXVuwREaU/xehxuCCsaHNihGcRRFqL4rSRPVA11kCFyjnSiCFFoDU1rhsogp4UbY
3AUxHkllYoQKvQvOKpJ29Uz2Tmgq1byC6chwPd3LmA1Zt5KeDc0Wurb0LdK+q9TaS8rj337Con4o
veYdrIgGtwnJAM6jnYOcH9/F8fvIyGVnQm7PGWDRraKL2HSwFZZY0w02hO8jLK4dJqNVpnuCq3qV
GbICrVDoZLn1CXmfANd/2v9LnNoHk7AuY6yaNDxdhxYQTlDjOnU+LI4HXMZEuTzp5nj5RmImuQQ6
mAV2E5yPOI96ZXl1X67Htyay+QFc0IECyOyFUVz2PGgkQMkCWFlA3n8mI8lOR1/MRBEmW5FY43Cw
C/7r4iQ4MSMBNPRpWO6NfZr7B5nUuvlvVC96keQlOlmdx4TuV57awTHRQQtKqCtyupOClFJFkyz0
qBD4x9Xs1Cm+cc6J9Y+0kRgCkeJjnkIRZtmks/55B7qOFUTzMpfqMHKpCJ7xv8GdzKsEBuGUusOD
1BRILVo9sNXAQCS/Otzb21/c7WNdY3ULaFPqGOK7DUdSzx945n8TUcDakZvM3vzdmzEjdrWXjCsD
CHGO017L8RSQYeGTYDOM2YhLWfaGWGbpOnsVEM9f0jF5ltiaDb7qbdJCH35XM+HQDvfhpZcowEdv
97OTaslGd89DLJhLx28uhujp6nEok6Ca/PnhdjhG0riaMqC8ZChwaVJ7HL4rAhuvXwQ5NxqLwln3
iUkC5afX0kCp6XPvpnee9x8tEGKHDUL2CQ/4YjhAT+m0CGgdFf6IOxJALocHa2jH6+pmeMjWfD/Q
jq9lV1xbbb6nrB4rT3boE3w91Cq2gFRFZSRVlfJ6dvgGvl6SqcirBMdlpQc1mC7+eDOhyapKegG3
dKjISYz0hpWD350gg3F900WY9czwAtR+0LlRGQCGHRdG+xTrg7kBTYvEcX1r5gFDHPN6nXl3DUpm
Xcu+3HNERM+J/s4aDuHTbrSKeK64yO5XNNh0RGgjVQgoSAQhAggKCWAng3w6CjE7LYZvlwsAop5o
qFR/+kWQ97QzjshPBF17OE+O4A5Xho7kEte3LOngP55HcvEE74qjN2WbKqw//2umGqu/9w6eLkJq
P9g3PKBU3Vs3unoh3JSJvOuxcpV/pPkRMsMI9B6dLq/f4OWry+6XFe/gRuoSncgmxJ9akFfCHWN2
L1gvaG6dWciz9Jx4tioBuoJx/+0wK9hJ/0QMc8G9zcUZaz5qJlv3dkckndsbpN9K07MkCl5FAH9f
6pH+rraPVjD4s0GGG6Qeq9qWIBpBGqv+b13aoTUgbqJ4X17M+j9DFx7gouGgsMK2iFY4nbhKeP/o
OxH2aaWk4BdMlW+FSfPxk/om+Ohg12u1UDOII2A+LZ/gOPUARKhkkIOsGUiTWNxoMO0ZuJ7lgTf6
5b2kYqLP2LFTT1ViJmKYdeyItZUJFYhzeQcpaQF2j45L0fu3R5pdAHrjFbCjN8cBQotwXH0O1y+E
faAlWWVbiiv1MCmb3v5B6qTNxcBZnHZb8yT6HqC4qY8JUEz96ZRNkwZc1+hntQVrd8ZBRTzbap8i
/tPxI2j+WBe+G8qbRDSs82wkHj4mciRMv4v6KySxABlyJ8q7R7YHObkbNcxs4U4GrzUSgMf95vO/
c0cnq8u2NUALkZ2hKCmdceT8Zi2EbrUd6drdBt8mdkmIUBZXOF6wqs4iiJR2TAsmK9O6qDvSHvPh
8Y2/BedxdYqk4fyZIGAXPFXqHDMVyU0HobgzJakGSqnw6hGTYvyPCJz/ZqN47R2IaszKAbOixKdK
E5xgm3FvnaZ1iTGXmSS0SkAlY+VdGAYMoSCkObq95fPNS0G6Q6WQ1lt40R8oAPBSjWHR8VBjsaEn
tudJcJqYt1x/e2foOA0McDapQiRsIKdVpzI2cvKxvUTDvhpNN8gmdqWDYdU8ONq8gR58corcZUPz
hNkE6UqykUKoTzR0zs2g/FvMezy5u+39XCoTq61PgyCp50yE8u7sTrMclFhX0AuLypWfev4gj0tH
g8gj22VOqkxYhLEvET5WJ2/Iuxi5QPqIBikVriz3s7OJozX6LVSWPU8+at9O1PFvTMjpMgupLqdR
wFNw1Dhp7q3NjiKyy5mXIww8KBFWLphhnuivMNstNu4rYf17mHzetEtOFjiAtj71vHcdu4krV4jU
7myLPSzj52kZzXFoulDr0T5QAzFsDH9bMAZN3qdk3wp3MfAnMgKhyqVRLziTgMM4UMZJ4eVgCP/W
k8kO+kv1VBH/myLfVRiHZ5Pf6OGR8Ts9uGJtn4edtURBA7Ra26DObjdVo/6adKDzrcqZtrYKO/G0
RtfzNXh7hFj0PuzqfIt/v3QRs0QL0RGYiW1M3LwGJEnYobC0htYbg9AK8nvupmIgzu/uRFuiUWf1
jfnwWcmy1Sz4oQROiQ5VzXJ8wY5Aa/BRAJneaKdNlV/CHBAA9xCNzktJkRaGZMI9rIrncjYrDmrg
NOQT3RqxyEYSL7ODflPUTXHf4h57cfbLXhcUhv25/OjdePHeJ22D7E/77s+IdBoTismpjUsmFB+Y
EIo7p0hw3JI4SDv731TMY5qcrMSlcGhslxKCCxG9rRoM+l0uKtvlTpf/P6EvahhLJuh9urgmVJ9J
cQV3wWEJhhuEertXmZFHBGzeROUPo7H8L/q1FlF1gJFY1G79pSdHaADXXp/tkg509zFDavsPHbug
3RkEPOeIgPxPR9cnNvkwxkrtJGytva3ecabWDNaCAi4hEwqMNTj5S0yvJ1a8csnbrWC9j+h6Uzea
kB9hXbF/I9xNJK9IvrC6Bxeg53Na0Lr1gMpSn/HZFKK7mJ3SAUHwLIPemQe61l/HuSkdytZi+Pgt
XNHbZdFiA2MhPlMafrt2LaJem0DJSuisEv/oSVnm+qSfRaxqLVuOUnC7iqHHCQ9aTAK3x+UepVXL
BZ3C0TsgJGuRamJNZEyl/ukgBTNc93/1bX07kmV5Y3S1XUJIfjR1groakXgiCT6XVf1xn9hL+Eu0
ctX5wukihvauc0LGotMbM68dscGoNNUIFTw1XCDDz+lMm/EQXfwzRV2I6hU+adnUOG1umptznbp/
y0++Cf8J/YL9u27pKkfEdqO0Z7c1poxLItTbNW/7fP6m5kgw5X9YMsmmuZRQ7DZQ2zY0ManIRq7/
K31xpv6wWBC6Ix8Lo2GcmHaDZzQv4rqyVrOQVkmTSm/W6oz6E/EXjrT1PVrzQorPGL1bAUUo6Npm
WnYo5qM8vLi9DVAMpVYUfhrN2ZLTwYEbnXVc8E+ENrvRAPEocdWktHpEVF4ufSP3KT8ntp337ZKL
tyINKOTlDdzkRgT7xfi4N9u8lDZJJvpxG+Wj/XSQNzwuEqi95GxkdXg7I1wf/wgXu08PFoPowCbr
iHLE76LzRcLYssxrVawj6auDNrJVWatps9YEh+0KvkIDlM38ebb56ZLRP0/GObj5jt9h5Me7Dy/Q
n+MCaxuqDvESPZlyCVGnfcfN8e3n+onmTT4lkrG5h9wAASvZw+fosnTp9nfdO50Pevh5HA5C2VH7
GuxtCmgw3xb0+75MkMQqKd2p0JxffftXY/runYG67iV0bXA0vzaO67uPJ7QSj2+CETm956TP9Wpp
hraoTDO5yfsQbPEGGAUPHNJG1ZEYhlR2SLVF8nyXcjijDyhoymXt+6E9qbSFULg33nSLMV72K655
M+fSe3IvkuwVW38Bq61PBetRp9B9qekkGHFHW/0PY5eB/XwDYNmuwDnmkUIUwquaHJEUd9DQ2+e3
AID6niLdzMX/7JyQESs9Pqh1VqwVx+b7ZVJm2DMbSVpXdVcNxYE/JmQoOBzVdurXHu2OnM1VkHjj
MacnPlaMNLvDG6ysyiolY9n3mq18zSyZLx0uWVirOuWXaY0dSZkB2K2CxOHelvOnrmdDN8qdSDQ6
4gCnGuD4mwJHNadCJSr8EIU/AxXWmGPEkMyQYzad9CpCNrqWm3tYpNha2Y8Z3Rgu+e2yjrJUM6fe
eT9LeBw0yf+5ZwT1nK47qcTvrxyysx7iaHXff6jA2sAH7OInjegxJKFWyUxX5lNBI1Xx43L05kDd
DlsQ11VlQbsei3vv1x67eXY8xTddMUZTmeACES7UpzkWAoU74BFE867Gb7qSQEz53F8KseX7+9i2
ruDx1Gt+JDbb4z1mdgoYKpTn4ZRP/ABHZGE7nnNoCU5h3X7uBSZDHPxhQ3E6hjpnslpd7azAR6b6
r7jaXDYlBqvh+MnSUlnUrhNEwro5UmbsxJZk0GY2Qy9xVeEDggrItLaCipD3mxthv+ZbSTrKZu7d
91Mvs9C+m+A4g11lHsW+ztoUVlSmgOkbJsSzh7X7uoL0R5xJ9cyW62I4IouAyEyg0QXpnMWS3eeu
6fRk5SCqgasFjw8m14xRP/1fBeMjRKJVgye9w+cHFUzLyPbN8pA1G3CBO2DKunIQUMrZMwcF1+m3
7pcBEmw3OaEcxCebe+B0jADsMGkYwQ35R4lE6tFFEMk3Qw/8aBSxB7HAJqIJrpyk4ZsYfx2XvUqV
s3UtTjhjpwI7WpnSFdsZ85yprnOSi41DRFaLzMlkv65B8HUtO3ZpYDy7vVAY2PvsHaA0RTed22dC
R6SgO7zTBhaorgaYwDDZOeHaI1V5jA22gUNzX87wC9BS04DKKb7bvHXZYSG3SpK1XKNAggKzSr74
wOWcA1IDIciDeQ0JSkoUSx0STvVHHciPFK1ObpYZRfEqneObAWyjYTasxzwA3siiN+HPEhCxNwtE
qoRreIyezE8pa4D2hDyqxYHOd4BLS4I7KkEw57cLzJcio7iywTyfAZaZsV7CkNkrArOWaVdqtKhD
bR+XdYgY/oJ0j+q14PcYr2Z+/IFalYxhwQ27qoqNXzd8IzSS5HWz79WyX3FaeTVilsYOaPGYCjJD
5BrzCNQl541R+ttAHbyzwya/jO1nVIVzwMUIjh3Kf1e2REIA+d8rHGTbSZUd+NvbLOBZ3uFVVYpB
gAt3l3Yfi9tOpkLwdiCwdX+/JeurRZk6Y35sbQ66RS2OhFyl14M9CE5+Wip/8KOlkcfi1FZ+C+Rw
TpskdWPKRbcrGfL9HFGu7PUPXuT3LrQWcK3uhciGcQMAvdNhrDQHmXfmIqJ8JFRqCfLGMdcDsbwk
scgMO7XqKh+TbKxXB/MzWaSNCTaVi3cLTkOnRBg/3t23CcfLFOiLE5Ad8SWSFfBFDvPBAXQEw4UZ
YwplwxbgwRksagD6/DaJQo8VtdjaxoqkLOsNCMpdOxSpKdZWOxqfiN+/seRMiKqjFexysHJ01DpK
1sjyNr7btS8oMPdVXvfPxtGGxiaXFY4wZ9aL2XGuFv1mnmy+X5J2ZeluzMToHp6UWq7tjcBquLP4
Oa4Mc9nv5Iac3oM76QkIy2EfWBJklY78c5cTdm6/8LyISFficPRUAjZMcxr6Lh6jCYtvziO3fOER
Zx8jbQA/2TPD4gmelEbZCTi6fUhoe3aHIA9mraWmUo6T3n51Z2zpWvsLnYOylh/W4GXS/O0TfEck
YT44vWyP3TbfQHhJMZHEehkVnqDC6wzIc/majyMNLzvLsehYLl/dr+UGwkqs54g98QNsoM6ZK9b/
qP1C+ziqjgAnAfPZ4xRUy8BrKKWbW2EPehTVsd0aYrH/WM+/YwrRHeATfCrpHkkyNsAeaHUTJuDq
VBbrHeHJybVeNMrSOk4mbkFtANqalKo6ORuwrkEiSY/zFvmM6rWCTZRYeLM11QtOA/TAMeTuoZAd
hACq1dm5+3UCtYOvKwhuXhr87/COnxVyA4btbjWFvWumMNNQZ7el2Luvs7ECbop/n44sSHR2NPvb
g4Xsvjm4MJ7gxLexJuRNkPrqybAnrE0gD6E5QclTc8/Tr9bEDDo6e/9NguA3tYoTz3iZlg8DStYZ
l4wCjuYfA5HVrJmY+v9/4YaoSWRA06E4BSMJYvrszbcSoQoL7B00kKfqr8Qj+rAYHDkofXjcmvvF
kIGUKlTSs0W2opPmAepeioKhmcbEy/vj8ajoOhY99CuAdEiBM+kxMb6GY2HV7hSe8ovL7oBmSnEt
grjalbi90IvZxh49PjPrZ7l2JGoydBS8m5fmyiK67qdKvgKr7ICrIalq0N1AcW9070DnYzsFL/8e
N+5fyZqwC4D+zGutEk3Jj8SBxWw9L+fvBgERk/xeX2trl+nYvBj831+1zytYOcx6GDdd5WaKPf/f
Mmhiig8aK/L+r/ErbHvmoaJSxFlEytMjRvy/H+CmUJN1fm3erQLNfgPAaabMTXzsEbU/CxfCujI2
RPBu94GbxMWKhjKoPpvlR/7Cvk2XojTy5G+Kr+01xT0/vA/7ElGrJmJCMSWZMhVh3RHb8VJzraqS
QNdAUfi1agVxgh+dYBzYg+K/2xwl4JM7maatJ3SIPeo1NyMy1v+1OUzt55fkAW3aXVzEszqSz66A
8VIzaThgP093GAqHRIBt6IysXwsf1DlDEDF7elFf6MRbwKir5PSjepWHft+nuH0vVsjEaxEYddqy
xb/2jgUZv2+b8SKNYiyNMmofeKaR0dyUl92xFz+lbsYSaCcx0E0Kk7wjtVSos46Xh3cQBguK3hQ2
XUk5NY2b9F94Aos8xxOigJQUBvrTldHu94FZb3psEGox8mtranPc5P98bSfkrOYkfXyrO43YK54C
ZyVfVZHFW2ONK047KSMtw0YP3Nml8zXVaqI/PaugOH/G94uGphsBF7HSDQvKrzQdvn/zjuCfzZpJ
lh8WOQ3dhSx5fcoLkj3j0UMjg1BRsef8miREqnnvqnCabSjd4WQTW8ikKS/a24gq6b4lOXIassyn
1h7XVyVejciEDAJb5Y6eElRX2Gd70hjTY73p/thITHsgYcj/wqxgoP7YsXqVn2lEmOCImSL+syMe
4vLe+PCS/NLqwKbcn+nRQLKJVgAc7R4TOI4UVGh+d8bisgSlEpUlLhr0CqMsl8v79ZOKSjkG3MDE
GqFx6rLnfry6HdVk0VWdSMQmMTAqYBc09asLbWCX/uyfbwxoP4MSrA0NGv4mg5t6Hkt8FobBPYZM
8g9l3w5BlNdHxL6vfS7YTFNI5vH/oUHVsIfAKTssCymXRZzGgxjul83MagtFBgZGmQDoos57imBJ
K4Skq7rKLXYmePRSL0wxj9njOmQJ+8V25KTPkkCHHzUwqqwK3EFqoOMo6XpjS6z4obFtMUU9EXbR
j5pVFCmc/ssosN/CTM8RsfEZDh0wj+/gM2DqnbD5IuWt1PKrpYzPc3N3RebejTN8DI206aLP16QY
qCNoHfcBKEx0O8pMkprpPEGGM2T8IVNYBWeERX71cOLDvZj7Le1euMF8kEdsfNOxwA6uB2Vbg7Oa
HitZmomcMA/eGUuZ5UO9mXYWm2jVRSnIDMEj+TPx8YW5NeaWJk5HUp/pfNLLD1/v2+sHMH3jWngR
N9PO96QWrAb8xjNFJd48FcvvnEAkPs7y9sTQ7cotcD1MPeQ6Fmn6p6IiPxXW8Bu7k9+yLEpHSE+J
8usbruBmTOkceYMUP/gGbDuHqUlTf1L19JVy4GQwvpuHmRwz2LbeUttOI0LElEJ9s6pWi7+AyoDJ
L2RZJKaWhVMZDG1Ciu6y7ssrlTtyjdjGeBM9nQElckUR1TXvnocjCekkTlRRyjeqf1mE9js92GQS
y/DJPewsLchef/VtYkogYiai4pEC/aaTw7riYBxWthE5UfQACSt0pKLG0lUZnxxVnbRwJF4cy8TR
4+EfkWAtbizHSxPzn4AARyRhqZnwKp0tjqfCoXSXUbdSnFVd4yW6O58egR3z/rOG+QVC4g+JS4vO
OjsS4FuTc8iT2fs8qhgKt9WxJKMi5H5DbWKTmuCMLei9eBi4NohcJpsQjOp4FkDBGzLCT51ugdGU
GPQXEq50jdko65WDbCmoaWl64FJGsXw9roUAja3hcbN3+765oMW9jTYoW3YiqUQ/ey4BApc/SAZl
8mufYltlqmHie6i5nTITM1sWfqGB78y8fxQlJKiJVU2rVJ5ogq6lrI4VVUTRjO1Lz/h1dGIVjbsz
eOj6RF7SARlgVl0IcOgxuJKpJzPZRTMCIOrhXvOS7v66h0fPTsARRuNnK1ZDoDMb6dD36uBQ86IL
3kR2uV7XGlDa15NfbwJ6euzmAKm0/yAS/+yCAfgQplrTfs70eI9xCRdAN6OdyJd4XqVz/Cq9Ou+v
BYm47/+FVabh7wpK3GQbBZHyvEUMfcm/5Swv2HdKBUz4xEuC2MI9EuzccMWhZ9pdx4gqlMB40S5N
3UHpxNgXcXsW07ZR8Q6tV0x/GylS/gWfWhijnr6TO/bY64xF12OVUX4eTKB85WSyO9i5YSeeBtAq
UTGSi4pR7ENLms0Auw8pVG/r6hF+BfBiW/7mUuUvYDa1xTNM+Ko6nuNRFz1JyyceLgbN7V1pqelZ
uRM6tsw7foAJoZOCwHO+1SsAuKhzjT3EU1B+Qm5la7P1tKwloJrzfHHeGgpgXUVzrETv2w3ziXwW
2PNNYBzgszp2Qy4mt8/pmyFWW+VyizP4p6Dxp3kW4vmZHh9viSXvWRSqnM33Xroip0Po/JyKhhju
J25ZuRbxTo4cs6q+Uw1pLB9SHt53oeP+BdpSLIyptinJQ9osNwRj/qrlIef9vFnFtxBGTaB8IhZB
ydcJlXiWK1P4qdrM4jgEnzwlliZ3K3xKXqDi0NbLMHK19v8H8E/QbuSgeE6zzjdPRMp66MmWll91
D4VWI1KlzBgJsxps/RwJgxrjMTdAPkuAjV/F4mW2JIgZvn5MCs0Pg4bEiXpoz8LCmK99+VFrKAvr
5HH99RfnF4IPMtgBSbTq7GkPKJobuvQDMlwUvKGDMdtNXEz4dkZLC6x8xUskVh8jjHCH+QmnZOYj
aa+HjUSnc7MPoMi6F5TX5wdvsDsRIalszF2AD1uI8LGnQVtnbpwkn8AY2i2KuvM+6L3XYHwl83dG
xPefMv5XZSTudMZUZaL/vx6+xzkibqKywoHKY/i5AB9u+jZw5Pi0t7beF7QNK/F9F1DpmKDBopYw
53Hql/3mnsjBsvcdRzfX9yvVlptnoNsFfRKPYBnOyHOGvyPbuEWDSK/En9gRypKU1yJZ7IO8iUeP
rn/WX8dXijGuRWwCkSdoHjNm5xMVbZhtbDiIaQXbcGC9P3j9+sLLck6TP4/xGHUrMyEOyFm5yKjK
TFaxAsYE7Yo4gVH1MnIG9RsxqeyV0MuVPSosJJjbcGE4y6Q2+3UuTT9z0/TP7dDpJvfkl9jr1mKR
7QdR+g1yvB+vXedOxDXY3Gj1Pktm9sUHA0ryVkzv/kBAQ7lV332Agzjhoesedpq2Xyfd1pumc6v6
ii5n6j0ii3PWtUdo3Gj2hgoOC9LFpW6pxTQSVyhVc+IS8LmMJACQRLhMUvbAy9UXZIuksRAvogj/
UQOevDQg3ML+CtrlN0V10BwOl3s4jnPRUfD4hizY5Nw1fyIX2UqoXuObWoRs9cJ2cgsRHwdJ8qOY
SknIXXEhJ+iaJp9Tjj06aVc3KC1DJgPQvVDxfNlbsekxbS6VgeYUaTazHmIfrPNMyb4bZlK03KUi
K1qULJCRJG2uLpV6JlS5VBAjTIlEtAq+W6v+kM7Sk7ev7oR/eQwB88vN5Gv/8bfpnK0rxe41YYk1
4DruPC/Q6h5UTmm3eMklVxBXHtFMM0p1gsLyzrqMgh23ozvpJhKDID4q003Lugx2afnYaGBJc9uY
BAMSIEYagSt/7c3NQyhsQ50gXGCTD+OVmiu3wHouyf5iNzLuuTRIFUwZBCqIZbyUZSAP2NwYg9aC
bosWrEFeCN0oXOQYCO957OzBj8K9q5UpRDMtbFv3UZDMftUSTtBaGg2XkQ3r0sfua6Khf6lkWv/6
v43+/D9TDOCDMjNJIxpaap0SkyZwuWf1P7PedQM5xZGEfc296lJRvrIurxbjf4gXHfIR2KXrTsLa
y+S2sE3bPb00NM0N32zuxEo8vqpZybSIQalpxJU5xccugvwjE42cPVJALaCRWL++SkHKEGbXO6/n
ZSJYD4uFHT0Myn0DPxDC3Pap7doLLkAkAYVqSuzWyvsE4d1RQ70dtrTJKnN1FqA+YxjmnZxvxd4/
8qkxC336pCHCWC/uKBPp4dWWTrOYiAC5nu5STPNMSpXoyt7H7cXKmC4esaCPQed0udKis9pdvsXJ
8qWy3s7LWx5jPyJf4QieIZP1Uu91QKzlg5vjI1Yo2ewFgxyp9vb2XMQc5N5vvkEjxdMQmoZmmc+Y
lK6uFfQp3wF3wzHrcIsmYVbuuNdxP7UOMK+UblIbgco0zekqgkI5wuRg/54AFiFmWmZbD3LCcXTn
VeNF4+QRsqtN9rdqY82qkHq9TuD1F5lCBMEr7DqHcr9Gwds0TJxSSqZyTuAeimQa3GXKorqKRH5V
n/Rzutu0ZJg1ub6Ihl83sh1Akdh1iMnF6VjCQTANVK3nZM1S00GhxaZ2G83zSX+SZbI6JNlpQyfb
NY+1jnt33OOXLOEKT1VGtmid+kXY+fkqGgUf7l1GW+fG3atgOBHvE+j8HESjUSYeMl4IG9kPDIz2
ePC+8aBFdHdTifcC0BRkOa1u2Kb7rbBJUFtVuAQSTQE+mY9ARWLP6BeIZpELpJI1/b9yCuFCvMW1
j53dmONO0kmRMPmdaNtgZsLNRvjk9n18Kr0yNQeYIs6HN0rqE9n2MyNpPb8zyjhoiVVgLaoVZsRw
Tb2sZvekJjpWQWsfs3t8DyTgUaWrNJQSprwLZ9+0kHX9l7p2e58oFwc3Mis6hpZHZmvcmMN0zT/z
qYBdWoKRecjmfxD/6qOfNIT4PHIRmrgDM+Mf0O9wUxFTXqFe7YE+c6y4zhHCE7qlXH/cxhNiSp7W
y20hteHBO/Ut81kG7XVct+34+RPF3hnThwoRrQLs0ZkN8uT+dX2x679zSfMutUj9vl4Efqgf4FVs
YF0FJ9z9OmmGqc4QkMeFRXKKacNyD9GYScPYnrlc/gF+ims8zmTlwuVOWpV14rtePozYTaKcJNQU
i1yUSldU3hj4/d3c0UIxfUkpKJt5QUDrdTNuWi6jv491dlWQ3ZSfW/PR+DlylyRyE6hUdF8PORnW
9ZmcP50Jl1R6A/3NB9pk8+4N0DsSxSsgbtclMeWLThosAy91g+SSVBy6DwgWs8zenilGCji3JVe1
5WM20vKonhpUKJXVEA+i1WUKc9YdGMgGiJTmVxM/SmwA3LtHhIkhkqUP6Ka4XhABM2eEI+XCdRP/
FZnh4ubVFYc/RGHYg5R0YnCspp5aLv3787t00BqPGn0XWzteMNx9yyw/4BQ3kdqrHpKpZ6z1LPYB
JOhI3KqOaK/huHz7+IpdPdJCT8+CpT0nDXmO3o8UT8QuvjOTj4GHptlvKWibWkG96IV+/yAulVgU
ihvskPqFWEKpoIlh4ykBjIQezX9HF0sjed4j03Mmyeri/Jo+j3+Mf4akgHmYlBiQbzn8TzSJY0rS
VkRFlDez/93pdXOPinK7DTqI0Rx2Ov7DKRI5KAqSsSHZWDrezS5v7nyiiPn7s29GMXcVP3fZWwwm
eYsCbwX0rfHYhc19VffrBuo19E/zlMTEO88N1wGFtwonaEteNaJLUsypEUjvSgxHs7Vl/InrZMoO
HcGHAw5FNomHFd+sLOvfUVovivHksjqxWR9vAxw3i6uk7/eabLRyHkYSs+syLjwzAUsk2c7/M+xj
ygxOBW+NXuiqlaQVhN9G2zS1WBtmcMQi/4LKRYFOHrIFEIg0zjEeMnfQaKUU1ymgy1ng2EdLHy91
0Hqr8dcElruLeSK34Id1oe6ICGo8cvMxNSug7Ir6Xu5okMB9DzpQXsUXXzVDeVv1Q0xvj9kGBNqt
rSdCi4u4NiCYudcOEaXMqr1YSUCL952jFLIuVDv1c6bFX/91dz+qc1WiXC5pLnqGNW2Bz7T1ZO8/
urgSUuWYIN/5x39A2GaJhLrh4cXa8TsFw4Y9agwqBiNrLZYPOxtuiw/BQYbjAFmjBI49W2xmyUzI
JD0hDLrp047Wh97sXenrG3VsiNaNe8E7qplkhOEUmyfuQlyB4ruK5fGy0JCWE+iOMkkAvr/fH9/L
axC1dFeFbRYmbs6PtXfIrmfbg5YXyUKymX+p+ARQrgcKtWWRCimaGGB/ZMGpHGhZJESvstPL3s/a
rSUMucQOeOnltj6xXniGmCiFeQb1nf/KNoXAABXnsVvqhmWlp4aSWp8bQHyGz0qX8unxSyytehU0
UWjZMI3ZSuXoa0NpUvzkwVM/74Tc2wYCS4X1aN+1+Kc8UdCUq77Rk9soAAuk99+xIfgZecJXEnJb
dP761qlv+dJiNLn4qpGSHlsBZf+Qpi3qyclm9F4bgHP+tTsug4UbH1jMlwtmY4h6JpZ/AAzSI+pi
WkbY1aM5Jvv569ol9GO4IavYwSlB5XkbCTFalB+yA+L/g9aorPv4lx/ae9BYggCteuacfEfgpqD/
JnFWk2jKBsWMonbpRdRSTGczEiF8cRov8TcNlJxeEHyzO+ubWydv71Eojgud3uK7lsJT4wS8jIMi
tc5ZJ4lK+EmEtfODm8ghyME1zNAmm6lza7G/bSNMLzbAFyI7HupeBsEH3PkFp8zVMrdravmaA1NS
zTSpO4q6CY0EhYicqctGs6UJRkKFOcZ9JE09LBLu1jhaSF+sXUZHPXqtgGoHmrZcv1l0tp6QbmTv
nOW+qJ/U1TIVANF3f9FcovHa+B1ScBS6i2yDdXXuvC9DeKAPL+3J1LWLqMKntzX9T2YDeg0nfRDj
4Mdv5K3LVcST7pMoCzfDg0SJt78WFfZdUEcuJMoJHskxNdClPNbQDKc0dYm6G4FIp2kwc77vbsFV
plKqiDUrTo+lBiOp/IHJKeBttwXDqkioQn6t1ylh+h8ZYjeAIQogjVnFrIuXIllcNj32iw9ByZ8a
YKovD7+T6P2bv8S9mi1WJcEt7rQYoFIfn69KK6Ir1MStu3uTd6cmg8LgW9E/Rb1/rmAPSExSElNJ
xJO/XWPhzOSHULmtxIvIopCmE5D6Irkb17OPCb1L+ZFE5CnXTf1/1k5+Oc6cMyszuC2ISz5Gv9xd
6KgYUbQS8uYhQnEr81sZ92gQVA/yCqgRT+JNklQI9EhpkQly6GvF4KnaaqvYYWZS6TXoKQ63z6g3
+NdyD5w/frnuTdgpxuknxW5/X81V6zcuxbdgsAvPNndGDkvX54QajIWqxko3spGuZaA412j1tui5
hIn/cABl3rFLF1m7zXoLVQ9qilo4uZwBxVBiEoXN+kW4h4NMbMzBrVht9NfhGNzhCdKhS2LU6vto
j8XGzQ9giAERLiqKJ8aOyMNxhgghZkG2ARXd2wJQMZuGGSm2ZiyAsOJ7gIcvDXORR9feCy0hCg4g
8gqENrzZXVu+QqJEu63EoWazMbluVBfAhTHpS6FkOLMNkJn4xSg96plCDdUaGKEJS0uQw9oNEduU
qvEYT5njCNSX02S6ETCGsk4v84n0XAMiuRJ7ZE4L0OhklRNVMtpLeSO3Inr49uMFLbZdX0rFFjuC
9D6pPUhy8+izKNjsD5x4IIU2osV/ORAyg0QAg9uXkeDYn8i2+6wS7cqxw33g1rxmHHuRyqBZRusB
7GggA5nouSziZ6FQrfL4lCuuBPCCHPzr3Uvvlk6T3QmyirN4ncwty51K18GXwgKUvYTV+UIKUs5C
ZQVXEU7Ksi46ficRp89dkO4pTvQRNoiJSamPNpYA0BR1yWCRdYu1gJGG87ufJ8hLhC6JxpHIddG/
StoHZSg9m9Z/ULhZ8GeIQ3HcS8tz+CTXtiP8F9k+UprtA/+zrFaYJxiVxJnUOsPEQT09h+MCaCyJ
johcly9mILSolZDK+O6lqlHyuU/WBKOWUYBSjuO1S9eK4FokXvliO7fFssN17yVZBha3WKM1MBR4
CFp1ufHqrZpI2oKZFj/zxSUOUOMp8UeA1WiZAhaCtP3FFo2uIpeQJatK7CDus9DV5lKCcvldwxAR
gm3uNARpAg0kn4LI/886K0N6m/tiIxaUTIWA475FV9HOGHpoOytDj6zvzatjJrYEn3e3A3veie21
lNyodiDNDVZdHzFjtvmI8K6k8Hu3XHNXhPAWvAB0Fde5eC3PagllVuwwBuecPANNVK+X7I7T4XaX
G76lWOsMAZ6zlR/LcUWagxmdrSl4tRLwdsYveiZWF8AAc+kNg4hbAhlpAw9E17tG9pnDU/2n3KTF
sit0t5qEY0qXczc5eh7QvOPh4tCdcYquynwhzfbdPk7L0kqzvo7JDVleevbR1afW6ZQvYk4vfOUw
fIXJr0LyUcJpsBtImEI18sHBB0p4sTFh/LpoXb/UvuMBucDAkMekwDgVwc2T+8c9W9tiRkVp9z5L
5VoLfQT2oIv9npLylwGCbRi7GGC2jtwZsRpefV2krnVplcqjB1vB5v1ZtOVLGLltQDkPuqrU3msU
LpWXiA2sm+Zfy2CSH9XfI/9VQMG9iWWvbruZH/eDjK/X1Jm0iM7qti9Yo8v+SakjuiISkRHznc1E
nymdcidWnaQQiIGrAA/VLfrMgOg+S3AWTt5u/UzlbKR4UcbzI2PLRKWOXH1q0a9YNHJH3u1ZCeef
XDXaAdWlQD7Hf6mUx/dW7ZMhjsMX/JDqcMTjbyBYPRK1f8FQT+QuuHXrzXvunKcwX83WR8g5A6wt
wE0UjeCXv1Zhr/iKnnGf7LuxQrQlMIoL5T9xdo8YS0YtoeQjhETaDwwu/mRe7RFN+uuQAFzFvVLF
B8v+26FXQlNcxXJZRhYyZrmkRyC/6VkIhLSaOYsAVTZ/bOykkdtKGXr3OeVSkZUzuUKfrgq+liCH
KRRVkFC2oPf2BUiKgqXsSVDGmmcjMgaiawDa4zQ6ldhmhGZP0D7DmFRbIUXsjDJkRhtrQkACHLHo
rfLz1PV7VvRCvNrBJVLUcHwq3Ubb16W5szEABk9v5V2nld4pXjewicMrXY+GV+ROpUjF/TU1zDoP
bawc2xTsnv2XSXgcyFWD6K2KkZ47SImeXkZTaToRGOGfgwaiHIrybfVZy5OlbQ3mBOVZHczJRxDz
i0P/w7o00dkXRWRQdfxl9ys6GKJi1EeHdjS4ZfdLuLDShDZmODakD/ZjsQIXcDmQNrB83zijVExl
Vvs/v0bmMoVm5b8NKQGNFX3v3ujmG6BFw7Oih46PnnnO/wOy/uO1AiaZCndaGkoHPWL+5QSijp1T
4MiueTGkzAyv5Ibl4E5zhDpL0joz+m0qDhiW/aZZfHYVPGpCzNcGaJ6DdaFLQGbixkgthZ2d3iaN
iI2Vtf3BspyON6PsoKBKox/dijxkAFwL76fVb/mFyhQ2pN6vJAtidHre2Hsu31WKocD2DyMtQxU8
iFVB2Ka0kI4Jz1CHORMtGtMZoOUI4WmR0YuDTvfPNbhrZszvK0uj6MLkhmFCco+H3G/MSAPCn0jh
A/PcxeOO/TYO+4uynickgDfDK7Ae0RJkUNEKJ3vg08CCJXwUfV/YWIdPxsRtB9CMpauxQAJ5jXXg
GZ4TrVKkhstSIWO/5TAJI/zNhgJgO9SfqcDAv53bZdGeARqnWds/W1lUwDl+XN+sJocMgE6Jk2+S
hIT0TOJzr5XvpfAy/yTjkclTVIYf6YKGwUpBfQJN5rp/i3s8m+4pcPKnGDHsKYLP52K3qbwaFO2A
o9p8MXYOZUvroZ+1IiEURLsREkFi6U/JQgzMRYuR72O3GMgyTON/dSN/vZGJYrfuUBnqxufZb3SC
fYAy3p6If1iliTkwK7j55VqqlBjs42WtpVR/21/qlmzFHN/IIZbmrA0UperV/Dd9ag+kQXlUTSzA
dxK7Y6bbHCUSckQSLy3tiQ6ulp60eex/MNf+vaR4aHTJUAxLLasJSqIYLfZAV5a51t91gmc4Y3QI
K0J6UeeJiemWO5J54pWf38pX/DstKD87co2udgKoMSOSXdnm9/tFjRsp4yRQewcFj2LPHYLAwowK
WwtIaNFjuYQg7ZSQq6AySsx7+CmtDMCgt8j9KNsyPvIffCE4Q+VaFZ0E0k1P0f1zatPfkrrpUsq5
c7ES/ML36Yl9uZVpnfA7g6+jbgydF6d7xo/fFBN6s5+JxGWaHba4SC+/Q1xIFi+LhmX0ImZbvDfx
REut77mHZlm+ZKZ+ADHCHBQ76F4A3bXPa6Br+iFHa75MNlhAFsr/0cYJdSCjaDpf4QpXciPdPYmS
nqiSjHUcqghremvSr8MDQ4jIH+Xsl5Jk1mPBE0huOQcKsocw/xTzpcQP9wgRfYndkZGwHwnkaZWz
2I86XSIPiOOY2CQB9XWTc9tKZ+l+AxhJMXCXoyhthnh7sTe4NXX3uAp7HzkCk2wjEnKCn/Z4eZ/N
gbnyFwlfUOdFJ7WkANSDgEPk8gJEeowrkn6fezgo6+5Z8dTTbWH4N1VzMorsAAM3y9OK1IImZRPg
g/4lXGoRhV/NwGHdiF03dqAH4a16O+Y4afPL/FIeMoX0szaQlBZYb15FGnKTe4qtUL+z3tjAPUEF
j5dpLtSNtxiziwwBYbNp6NN5yRUCY6hHC1J3QMIysgr1dl1+40jrgo+jTQwUfMg7OLDCqR3YrLUz
AV1sy1UpYzv3OQr32FsNPZU+I86GmLFE7yMWt/OTReE3qOJY1/AJxkZH+DoVC+pU1oT9G8OiaZ6p
kramLKpszW3tqkKnY4ZmMvPWd5hh2g7sZqDgPCCWp+uTetmFZrc1pU0XLbyFJvfZ+uIPRZs0GBZM
uj2Cb2LIztqNdOHje9OpcHFiYCh8vlv8BtP2g1k0ECDLGTmt3OEFTjtIPOiB8ajwfheA3YWYeNoN
WJLhfTgVwrKJP6fK9QymoQ/HwG4lEeiLwM2/MloEqa/WiByLAexxU1pvLJNVmy4l1kL0UJXFVGZe
/0Ihi6OvfzhuiMWkvQWH81WoHfPHV9ztw9KModvkHPCsf0dQwLKzO4+JopLDku2x9gUyzuwIEF/K
t8Y0hD41M5GwvGBQdm4WoZch6bdHLz0w8267kTcHdsasQboXaNyLv5241BP6nhX4CZSIqtoeZJeU
fqlk+tFcKAJNA6qyt+SzE3CLdhNCQfw+wvxGTPlLuAS6jufewtFyC5ND4tP9Ub7EAbtAfa/ykzwc
7MCZdqzTrhbD68fzQ73bB+sOw9w14znArFmMwtgrZc97zIxAWO9qTEosLhFQRqcEm6PgwltK2JTX
vyTfpyqwFhgm6DwoDg7YL6qq3UAZ2muTor30dVoRoT2IYsPZxTWLbu6KGySAWxP9UyshwFPTZWwX
SlXKYsWJSeEnsiPpFFzqPYEIy2ZkedgaZTAG5637Sc6HZiQlkl9Y2aDthtv+2X7PpQVVm5T/typ9
ItPeiBcbvTIHC+pZ27n0v279d4uiP1YppZiINHGSKR0Imc1qaCpfaJGvzA089FSY21P3pwOFm2qi
IRDvcWaQluZEMDaQb+kx9whI+XrIGJ2cgjadBs5s7rD2BpGSeHm3KEChtBK0LLTTzxHEgJEkm4+x
kvXPTTVdSajm3wUDQbyYmcqsUwNJelfU1xJmdESSDedU3CTJxzX7yw7SZWtrp4G+XxRP+vq6Oe8S
NYq6kTMDwrrJ5KEGN6DZzb/HDu3erYBxiS03ZhwywJOGVRUwL9LxFpbe9vwSOSgxSNPyW/Ha07tp
pFs4hC2KGIHyx90ylIAoY0CvJqFa624BQI8iSVlvU4xGtcrosZwNS7QI6PtnRJ2HSiFjxhjLLZTK
uOd2RH1zeoE+ch9MIavD3y1wBKlaFFEpmJZ8ZWnFSkz4Cn0FrOchqLLPBWYVx+4At8gV0qnr4jOi
7Hqdu0teuo8AHOPVtsf8Y+/aSTgbqwXhQ38A6bLztxXbE9B1pv7VXiytLEOwkJwFFkdnWCjfWSup
KHGu/D3ikFDQ/H8VfQx+IA3hPgeBa7zHBhikl6aDLsvqz3EaUKED0wXi4YTmy2atX7fInUBGmQS+
e4GViyMFFot8k/ei91mdBr5B0EdymVA4tgwVTvR2a9AqnS4G29m7ufF8d0XHEUAAnmBSFezsCjx9
wvPSQnE1WquwkXEDIElhfrTfVsNwIpZhMjUAhImWzmggJAOnoFtM6uaLgfpOu/cAfB09Hy1SWuPZ
iYm3zw08msELklOPLLwOPilGjs2OCHFvBFw3noeQ/fnl4stKri0NVwHcM2WSp3Sm3m9ow13Ni9mM
P5fWX+9mo2qCaRjD6pR4um7o9F9S2QlJF3ygNgf8IPawtbPFrFwL3yRHIk3hZkGKxa4ALtKzCPwq
72ErmezcJoNdQoabOxl56Mbi3tFgxj2x6sYFmXVRTRha61q6ZBple4r/h3T+88MmC2LUkrlGVh5x
I0sb/yE9zAKOKGbf4yHEDKF3ZeVOYFZX/ihZV2AvZErR7F2smNETANinIxQ04auAuLeBGCvxIDxn
VOA45yMhMKoqFZBgWPXkwJrvMpJsdzV/H284nlr7bYp7AJTLYeZOuRaVwBM5lxogGLNa7p3vHBbu
3UQPey5rlYYLjbYGLJj7AGcn2CfQffwZUSV0ZaS1Cmlj/3hFamWF85XhOMdgNiq+dhVe1vxlErIG
BO19NvHPWRm9NYkqq6d9o5fKE/kZBf5MDDHznjgcqFq/D2WSzUKUK01PyY0nkLbbKtFavk6Vkdb7
h1XU7yCeoDfJz5GYyVvTZseKPpQwak1Dsil/0rZ59V3T1uVmQJBBHnvZkQFHZ21H6fJWVn01/CYU
dZV1OSb2lwZPFeb0GZlHdTpvfBiPuJkrXR16yFAlqhp/mqitO8FuMVX3WNECOA3bWohSebuuO5iA
mOnvI4QYqoWvl+oPAfTPySfC1Oeaj9TsC130wuwG2/WamPZt0JgM/lLvjGHT8oJ3Mt+cG82DsDtd
cI+1fL7Ka3O1t7smNhmbTb000bHZWNXReMuXSX4w+/cUTSIKWuj5lAtMI65/82wwlL2WsCcEEtLv
J9GkVDb3zMraL2Dos2cMmVSLKSKjT/gdDKb0JYF0Qfq3X5tUD1wJ5CDzcI+Y7EE1QM9wbYyGfdu5
Y6TYekdcf0fon4iuu6Nj5G7GSAjPNKb7BLdl5i2pCRGiGyNDyWjSXhd4NPVrLAkBKlx7FxgCmfTa
J+rrCSeqkltlQeFzW5A22VJ72oORe+XwIHYr+rJUM1xuegi8fE3Xj3jqSF3200yDiJ/lBLTSYw9T
8lzMNg22r8cSRLnLCcc9orJxorkarUE+7dJbHfdivT1zxGCVmwwZDp9AbqQwPoWx+hTkQQx1Bh36
CWpJVxv1v3ROsn2VVfwO17NPJfCG+P7UUTrvDEjgLE4ydQCq4e1qw5De6Y3+O4AYWEF7IZWu6Ugn
iPjY2+CgqAuFJ5WdTPKhEZOq88LWRYzbVrk80aXpGsOmmmpXEI7/DJYDSf3VDJGDLZNjsot9Nqpa
x00AsIf/NiJtQFEFs4RY2q5o0j4IetItUj2Uod4thYp+fdhM9NV7wOYVQaxbC6zx0AYdPcqMWvD9
Ssb1FGgp49ysf8S+j1p+3SwoqLkmKfYZlcOUTK2nFd2WuNYnNYU6iF5Pa9W/2Z3ZXVEWTie8Dqx/
1NgDhtHzWD1+OYnuWED/SUFKtw0mV3jc21Q9LV2o+090UNf2sILDRlPYr12TQgZ6mZyjbNmeGgz7
yGY3y7WJI7r8IhK/XfI6Rejh8YzewMBvrSZH+EFW7ibEXwkQg4ax0nqcY2EhMiZOpy9SebWIAiul
CiIPALKYUZiNd8biMn9JDEosei8REzatMcqond7uHRRVH2RjMzsuX3ic4UCpwgRNY8FNAfFp11HL
ipuElXj6lcEYZCXZO28mp9jjYtkP+RHtB6bEmlFInSpsmv27x44AA4EkT2s8bVgUyP1hj6JDDgDD
Hvq0/bwQXqH06TjMSM9AZ3Cmfutxe60xzlfBp7ihlSBUYB4WAq4ZSn3ALpVjvHb3utPpI/eMDJXL
SJHd0EPORBXFIJUGBhoWgTy9xfU4kcvI1aepLaWWwxHx5obekIGQZ2SOWRLNtoz7YCewpqKMyR/L
i8M3Uc63aeGGwkUemn7CGRtxIcepk6h5cSpNC/BrDvQtV/2tHSwVzyHGKDe6sZL7NR8hiC2S5mha
OjPlKPOe28rBHBp1cMfa6l5LCRI8Np5Hi+yyy205a1pHAcj0s1JjG65oTlUUYi25pEUWzTVo4QUb
BX0veNpT36FXA0vWP8FyeO9evvN+UBYYYk3EEsIgiC4JFFt3NkoUAXWk8UN9y6KYJsoh7tH/lrcr
yQQ01AEjyOJH4dOys8ocbvBqkSt0NxotkTCXfv5ILyfun41KHF9wVFCQ72bpi5XJJsz64YyhwpRh
JPocfQI+ySdMawTYyC615av7wwSU9jhpxpm0Ls8gmQelJgtLsCvZx8EWeIEKJfl3OToTN4dKtP6E
vvU7LzMq0S3qxJRbwBpBf6XtJzOoXylmNruwJcqQ+baNi/sVbr4S4hs++TvW0sOrDHwwmO1ttFbv
wqe+qB4pxuHPtFZOjDY9pdGBGdKh/oH1iToteH5p5UCB3MdPBvvQ5uLQ2ZtwJTIgps8nsm2MuiyA
xIOkMY+un3t6HmDPP+/Ry/yYQmzkxvckyYSNCXn3nwqPw4ShWnhXPAOsCMk+tybNYb7oT1pL1/XE
hyD8svxhjetR/79elORfWGYX0fLfwMFeDyZ0nj8iMwucEpNj3yYEwVqhL76JlAqL3CKl+dYJneVU
+UNOL1OLKRRc1CVFsXQyhemoOnWlpNkPUVBWAQtv/gLNHO/4Dq4wDiByL/2JZ0ngkrKh9qjd3AHd
C5ygMx2Z4HEiFDqGUt5+T5/HBfFST/glIS7ryWsbT7Dgoaygpa6KdQX4ZNz3eDl6RWQ/rDX5BD30
AoJOwiop3cwgTVBzF/6waOP/Nb15fmRWAiFgbf96po7GEwPyIFDaYtomtU//fqVp5FRaA2XZTm7K
KK0yF7SFfSQpeS0QypcWUrmNuwQptk4PLPJNiTcl3aMb3barfOs40RqMxNyNkrh38o/2+lbOArQ5
IrPh23eEkBEW6E3OUTRlqKyUbzbBBrHruT7Lz0F5xYbsia4BXbk8xot5XPPXZDfDUVo0f98KcXWO
J9WBVhdfc4auLohzYXxk4r8VwTmI0uY1iDpKMZfvNz9oyGXPwpelMS7YT27TDIzvK03AB1yfNDUd
zEzy3EPcmMiDXxpT7HalD2xoRHeZTGNetwr6gzEmh6Y9+7GMF5hxG+F61mLlfpD46xoPKylCQ8k3
iis9K5cLKaLS0vi9LVjqVSDj/KPqe/b5dlzMIzbgx9PxiWi7yt6JebempFXo/caWIl4PcMXGBCyk
h9ampNNnve6CRUuBPxXk6rgml+5unysGMOxKvlruytPzhr1py1dZmGnXkCWsoRgD0YcZf3pgg22P
rxkBLeiy6977TEn16yoBgmNqCsSSTnY21O2FT+DAdZ5bFZ0tDIMti2jqNdgI8hRB9DB2Y9L5oQlF
Da4l51CRG4TXslAj4LU/5pmpHUCzxJ6Ee2jgggVciYM3+XietLj415EwXBm9nmKth525CNM40FJc
N9K3cBo9y5X1MIi/Dtp2TyyM+H0JLB248KT9p8ocayBnh/i1Xu8RwhRn3nkqabVbEDTCBrHupNtB
1XXaXuqDQ4ehKMYG1HUuP6f+s23EAeBijPC/0xpjqVMq3NTnK9eCfYGLQJ3mBxCcdrIsU3iH0fwW
GcKUje33VPbhtWRWWaEB3s1gfj0nc+Vvu8H/YXd98Pd88WutelHQXgVogT3dPUHPzlBStR/uhWXs
z9F//cB8Q0BH9j2NFDA+wiPPckObECWSz3XuvYZ3xNzLoMORw6lPJbK4rn53h7rVDPDQO6wKEYMN
iwVuQMbXPhSuwVwuYJM9rHqbvls1uwZBEziVnlHod4gz+8gLN7fzq2V0iMec7pxz1mr07aciv8iZ
/Ap0OCJDvX+tHN3vABQCPTD4EXXPNGmX61NO/0w9xMbRZfmK8GDfNo8HARH4c/Db3r2Evm3g1nxI
dX6KZqVwkhuAKarFtey+UDrq/tqnYrQj1v3noCxNzSUlWw7LSnQyWZSqcKHOB9VJIj+VUGj8tW5Y
q53z2CbAyCinsBX3O65je7+rtUa298YK9eg0OVrTWov475phzXVp7wB5BKHdrNZMBASPdKHJMJ2f
n6ARE2tQj+Y3JDdO6zk/KG2IfGWqUfcQnk3u/TnCy2KtdpZzMwxvBv2nNvuFVn4eeXKR5XqaUaOf
rQBg5DU9qT0elNwPevCcT40q4UxAjHoXA0IVo9N1RVO0h8OeOlpsNiaf5TqbyKwp7T6H4fKoArZf
mW4ok0msR4/YURpt7Ek0DqWbRedt8yIV2zFiRh1Am6UuaYxVJ6FnXIgApAjVJHwv/5EAK9lSoZKN
ADdgPD8DulYC7GyRvByiaNEVpMRaL7Y5bppxgJ5U9FOdKF7Nxk8jzOSSdjqNi9igSIcU+ebFaZrG
vHJ21D9y5pqX2UVpZGO3O+sAf6VjMTccWZd/VqvMgDuth/wElayUTqcjRgPabNmLFDQHKONvQfAz
Jane/DaShyzj35s7YI1gZMTwwwtVxmFXm2A+ykg990od5iZ/50k6aOTpJWegTY6IC/g5IzmOyZAg
/KHP3M8240ZqBQDOosHyH1O+7x+0Fz2h+1HOjlOhUhce09IjJYNSdvFMWvBe+LWHEwhOhNF7ee9N
qHd150A9ED9+7dvjMWFcXboCBR2v6Wi4dcazIe2HvRY4Vh4DlBLWDxX2Jug6Vog3Mhbmei7lC7H+
b2HLJeERcEGYioJJ8wdH/Gay22O6o6e9yEILapvhK9cXuRDKUZ2qLc8goeKNug90vzQM1D+4yHrE
NRX0OaWkkQ+/kEv71oArIgqdJQYaUgib2vGcH1ADWdhUblo/hEqX34jJ4EGINK8idcxdkSSmLRcv
fnVNRiLAUG3bAA2KFv8StOms4ACQiDznpfWL6GlRWJPDblY/aiMWD+8GpIb5hnRzroV+uZTPHSY8
kDvJ9fbF9xp9dJQMv6GGi8CCBqI9NWzuP80Q+JVGXqbvRnY2EtbT0pSjKq4ygbcqQdBGiB01J3WK
LDWyw/1CKT783ihZN2SQqqTC6xLFJYHmxPn76fe7OYPYBRaoj4ay+UjwYKCRjP3jrO4Nx4BhIj54
xszzpLOdYACjsbajuiR2kJG1lIR9Lob2d0QmFZ29lhnesAN64wX4Xwv/izySHzBaHhUrKm99Xuex
GZPrDKthIu7CsBXllELEgYcZcWLjSEukYQhQEv/J40I57cZd622gjauiNoITsT7tsXpYUzwHk6ik
T8Lsdcp3bGk8xYcWT00oG/t0jURhZmfdKkekgjtLY0iLYazAe517ppNYMNZeJgvY+IGZMcmUIM3m
wPhZ47M/hPGuO6Jfu61mUYTtwgfzL7xhIB6QUP+rd6buWj7ZLSk+t05HPtNLXrhPKPN8Cu38wOSq
oh5Znbb8sGenG4CM1grzFQOUJtNlOexe5eaw0hcFh3yhvN71EgzKEYo2Iuc+WkRQPyOEVxEWjNNk
oDa/wZK30uygXQb1lCOnFv+/V9XNL4IcjIYFhCm9FwxusqsciDFrYkJ6DWpbSN7FJevPP4oPFjYo
o2wAg25vFX9mu5H4KVmnbUz2gmSXcDcQplEVab//eOytl8Lp8nHwGoPjp7tQtOvFE9Qy7AkbhtkP
59294YIqMsiq7/CpIWCPhuL56B2BUNW0RM2pE+NDx7Yg7EOaCsp2e3VKvjv7SObdH1L1/n8WEzjw
iwFlLHZfcO6exspH1xC9SJz0zzeb3ZL4NrpcR2MgifQL+T4AtTeFSFcbEnhicHeInlK2Y+ZtL1En
pNDA2kEkIRI6+lahPaAXf7uAGc2kX9sSUuYxqeO1PIXTdNikGtIXosZsy8b2TYTJfHf2tKMEJVJX
CMIJ1sLDFuQT+r/fjQPq42qqmWZd1B7RPzLExls6KaOUK8YrFrGbXAYKebEJ5HgiUHQMADqMDHNf
CNIG0q2DZkyxgDi4dUvzEjp04cmLFpnku6fpGeFSSy8t9mu0dTdQyJFC6MtWBiW9/05O7Fqg9LSW
7lDjs2MJsIrd0ni161oPa1WmhkMHL9yjFnAZDD8AzFN+rnzHWOqnZMMmXBk9d2lhCwzBl3UJ/NW+
AqkMJckqFgovNCEaeleWxa3BfEWiEAkpl7vdpeq4uwqmKboAai0xAqM+moyR1m46S3ZmT9aSIq/H
f6PyM5wwoTrfhpzqaf6l5Vi8+kquZnlTI8Am3FzOLIoJHflOxN4uVspZJiMkubPkuVHkRfn3IoJ+
igTsalQKCf81XUbXT5EWG8wWqnkfFR15d2ggWPfhTtM1e6TG/U4fmN8Njpf8iy/Sa+vDHB2HKr2V
JR9TlywtjM76OeB5ciGaiecjy8VPPOH6GnjTzDtXfT3QrWAUA97UCbEcalnWqbtXsSdsIyc6ti4q
FggkuhoYXmk3iiRj2ycJMnkykcstOc5NBtidnI2peaPCxUjQwFWDKy/ArnhIEdkf5AzQZTPHe37g
5293DPH2C/e9MC0kwUYqwz76RK+xxzbK2lxS8VeljB1jCjUKS6S8xYI4rbTojH5QKZF891s6jdGm
aXrB+Si8lPeV7hSB5fQYiTlJNT/XGnB03Mcjig20V50UazxX27NHZXihgTFToz8LiZ32dtGr9iOY
WIBhFyqzAI+n159Y6WFFQOuNGC7bfBeV8jYjnRPPA0po8msJ2xzHz/HVbrXQqbCgWMqVfkaEHJjH
lwRg6nh7V+UWHxDBO4aV/NEEEfHCgpzwIuap50FQZwsOKQQgb3GAYNsBOnj5q7pPjZgAH1tx3Rtu
V9JrZJkxLlt3ZgK6nmX1nB+T+wx3Lh/2hhI0gWjBB9lKiupOKHkQUkvX0FosjbwIAVEcbmWvF8zR
/+9HQ/yHq4Kg4u7yro5o3YqpNzlsApLLaLT188T9TtcMpImIbDMVohWer/wJxKSIlS7i22UnOLe2
2sbXiP4hSmtJ6Nvk4HV+2wcJmMRalJ8DJA6CakVa8qelDZG2RUXje9bp/eWHdyzgJjVC6MZFVsmQ
WmsDB89jE5zspeekJumPIJ3cpixd2dq11mYnibznE62kpcoZ+sLjO8+QW6dIoScQGvTA5uZo30V2
72vW7c1CIiaIA2fusOA4uul5eFqr/cyTYM6s99TNS8Dklnh0xAXE6XouUnJfTYOEW1q6wi7pLUD2
De8vypDP3HzGX73FyeGQKkGfZ7CBdZIS7++5XrRItBQp7yMQ8FhY9oQt6j6tjJNKwFuQCWLRf7uq
mNmnKSeleJPeri+zefsG+SjHodNWaZ1+z11WpvwnGXE1O0L8Xj8+lr7NwSQCTZXndRWGa01mZ9Om
squUxCyW4k2sMrC/8cxewTbeAUwWzW0+tYkMBnv3dWZEIfpbvvfydKruRjfHJWYXLntjKxavDBtM
TN5huPOGw69bOZPCXpmJgvnL1czObWGGVgGcHwlb7r4rUE22mktV4/YEPERXRWewysRsspVr/lU0
INxJ7HfXoZ7b4+sYNHNRd2q325ihK8IcxNCuMowwbprGd6OpTXLLQTuIwYXZ1szPDI8BGJMUfNyx
+euPA91CNgE9nrrJob0iF1KNRTx8tjNu/PaXWSN86oem4RoXVeBk3vbfz2v/2tdmz9d0pVK3HSM4
zHK2zW4MswUpBlzZxrFiqHfR39wUG7JopTTLhVFj+KxK+/RYTI/ccwFj1xgYEQ3GMFZ9XO+SeU26
/WgQT+litYwkwiUHM3Mwu6JcA7m0Gh1xMPQInYe1NeCE8bYE87SsC47Cv9JjwILt/dCaXiWScgJX
OZO/HW0ge8j+ksCqdmomloH/jAseW1SP44a/w776LUFA71f60K0QriD1mDw8sR2Qe7UjQozf0cdK
NeWShTuXXcV6hVg1fRAbaz5cyr4HrsSztzJYdF0Ekd7D7kQYR0hNLe91CqeWBjLyp72umK/rLFUP
gBoIfa6sq1UgtIKgxq15MikXeekQKJdTKpTf4j466EW4ZPsH/kFY/7V1Hwe9jeb2rw9X7wOeMD8Y
J17UoulxEgqrpknhfHWl/f+NyxP5sNOlQc+Lu/TZytSCIDi2Q6KGZxcf0Reja/4n/EhSO139kurO
bjsEM4XF9QynODcOtD2BApJK9sKAd7Wuuq+YMwJMVOl/sgQh1uhG2Mfev4HO5UWBZSfz3is4lVOk
NVPpnYm3D/dshCOLYPXt9hJms8TH8rXrM7A10RM/YNh1L5jDNg/lli83gp05M+HqZR5+mtzxnicW
430TYf7e3+UFvU7b6hqRCXn5SCG7BoPJSs6DCZFav2ECUbb2I0M56fnEi4DmCD5toBvQmAhsQRsi
JvmDPW9dKHAzYpfQu7NFIDrWBchrE+b9zjf4sNRreGG1sUHEOa/Ajy0h7zFthP8sePfzvfhi+A6n
e9y6XXHUCihYcJfAVUY7coxInb3fjy2nNQvyhVbbb4GfrPwdnWQkcaPDF/f05fHpKyUGONp//vNu
EtbjMoR6qdvtCPbAl1i9YE1xrUlNMIIofPdCFecfzhBwEKQh5Sbx71f31qtRxkncVCzR9t3jf4Eq
UV+/yaIXh3A07w8Qjj+t5OxKqB+q/d9eWN/N2lbOoAwc5mgaaz4YaUqjI9VSdNeLek7U7SjjQExW
XgJS9E3RY+PXqSiYEUKnVgkmLJJXviAAP0vPi+RDEt0Uy2pBjxw0YEnCSGQtNgiUl6JfV/UtS9Tc
Pmfr8/m2lj1h8sjAUAAq1SB6uLob1w/NmF/wPdxZ3eo/l8xB3aAtYXxvru7aJjuI97Tyg9RA+6yC
wtf99yMVajUJQhdK+ejJNPPQ74iEll2k3gpwltqdc1oAu82CGkx44B0H9f6imAc2VLJ7Fo1PsGHA
yuDwTS2EPXgoAFulrUTXgnuowYwH+yqdrGiTHhXUkF/rJo953fdh4ABRCC0+AwdTD3irMKxLMFCS
G/1v4LYV4f8y0bhcj6JOnHt4ec0NCLdpNfjoyQUpDK/ZqFHRkkcyRPnO3WXCaTno7dh4XHiivEKE
kcxQcRlqIk4tZtzJPUDWxsqwjhQfdjJM4aQ4Sx9gSzJduD6E3G9sqeHG7PtRvJ7It5Q7E5M++QJd
TbulgSN3YYmd4pQsoaIzMuyfsmKGqOvKLbGOIuXOOHUvbk3acx5aT838rlQXKQQ83IDTk2rg7dqw
5ExYLh9bK/aKkFJC1iTQ12SrXSRZg9JCxlQcKpACEro5BDgfgEP3JDenHlJpbcBmEw1WH98/f9Kr
vSISgdnxfFVKmHdazbV5tNFtZcjbKagibFKG/DLfARED6842Imxk3oYEOo3tuXB9zydCZfjd2lxw
L7CZh53bb8V+uzTohiJT0wwBpx2mpn7LfPd8YLESFA4a7c/AtOJ9wKgMM68WGhYFK3PP5Mm9CBmu
nqS+bV9q+I6Z7y9gycoFDyF8x+IK3/I6EBlfrWDyCOro6G9LjPbMWhgVk0kCivYgv1XN1Ps/iv0Y
ABsbi287GBNKQVGT1671Ri+/tPp1rYGq26RcA/8vnvSAEjkgFzjsFaI3q1qX9UKJ1fcSub9O3YMx
gemyw5omsBihiduoretsUTya5+G5QNWOOzFEeZE6PegEAB2g1NvOsB9m90M0XD82uzaYmuw2X3U4
UC6/eB8M19kobwr8/NXT/2x9jFN2NJYWSiIU9ySfcgsNMpz9K5Vx9o5iABhvgEKMQXRxzxVyTZOu
D23rEqCfned0kXEBqxaMEh4yxhuucNwE5EYuTF6lVqLnhOkyCK5L8Z4I/JTofXakO12m9QwEqDiN
ctVzISYjMZL1SXLUUStHnKt/lomiZONKsTXUpghYYJoA6zCX7A4YK6YMDq/MfYuLt8zwZF2MrkQs
uVQyOw0GV4hcW4gEXXNklHk4llmB62L/JiMBMk+zQUltRHCFULU/PJYVDVYMFUe/VHv13dhFf7A3
ohUP1pDdvW6PtLvCjNxQNeQOYM4ZbRZUG/YQZTLeRMIgxXkFGUrXbQ1PjW7YC0GblF3LEiAEHeH5
NLRk29x3e4iPForC6XVfRw3avjxtPwR7C4f12BmejAjij54rD32SrhDsBldK6lUQPI/D1SFp56ZO
mM+r7+uqkN2nZpO+2Jq5lvpiSzacNqpX/yfB3ZrRdU9ifz7lLzkIIC3teBidLpaJQb59g6iayqa+
WZ7uIP8PNk7Xpaa3c77SDack8V6EcUBmceAE4U9sRZamUT78zC9YsSUwg+QNnEF3podxOsmoz4qv
2bj4pwdDMEYMndCIs8AOwWOOcFVDCR+m0nauPg6k0DOCY2tbd2cwlM4OcCYZze3OrJrtFUPlJPMl
KUGN4vNPquwAMW2HuizvA0JxpT5FdyXvA8vybBjVVdLv7IuhNZVWKL24gRJEachPMmOK3b7sS7dH
HiYemH5q/CZ6IGns+8jiKFDWn+YWmBcDfSFsJXfX+eLgeIHXh11FBqHM0qVYw3GhhYuRQo1x5qEo
Z1LHO183ONaw3LXRPqw/T9WPcMOS/fW9qRAMZPI9kRrYhtvbKqy7KUuCdGebWcSNtaAJm0tLPJC8
fwKgBta/mqsPqLdmLn66gzoYKtEbsLb0DeKq+Ze02bxWKarAUT+A6fbCLKto0X0ir3+3lVXFUxAO
8lKuOJCQRUjT3hgHFNN++2Nbq4AngeM1qCB093xQwKSACApVkLB8puHa/aViFbZS6xyRUefgH6mF
a0YNkqu/4oaoVywtE2uWyoMVCsM4i6MYUaX+DlENcd8qT7/M0yHZbtEbxy00VzvHRFw2J81Iw0oR
VmCzHq6vr2wJvaM2GGF7b9zCy5vXAEhZbjGUCdHzcWitv3IqZTr0SS6F3shumAQu8hSKOjpkyXOf
Hmwt6nRlivMvVvQgSk8/5wqJy3ldVBNpylNz8qLse+sIr/X12bPckME8eH4l1JkSc+oYfL2RVkyg
Jbzwbu/CtSI3xBNCfJVPU+o9IklIVepfloK2NZSb0BtRV2G8590QwLNbm5rEu+eM1P8qcFnSZ5tp
HpleJ+yG9O/GqQB/MLBqTQUGDdFAcPzM9zI8iIhNEX4HW1mRyaInSSHcYP1erUG+aKJi6hnz+gZQ
WN/PSHi3XDEuxsPeSdVTqyeY9WDlNxpZm+Idvap8XpoKsomVDoMtTZnkXKv9M6S5fE2j9fXxbGlp
PCP5HZkKKUDE01ZTSJBS8kSz2gBm9gJxtx4sJHAn8iN4atpJJOx6olhFFIPYXa9WIDR/tMxSOMzZ
WIbs1yiKkXz4IG/dm74swGR1U+GqYwB3ILTY/qpOR9/Op6rxDWYmjDegU53RGpyR8usUdAtZamMq
x1YpoZoDkoa3kS8UIGDueXjh0HULCSiAhDsli9jWXzAwSYVcRR6j2M2hWCYCe/YbZd0lhfdVJF5P
uUNRt7so/iZSGQU/HXNadh8zbFKPSo85+4gdC14d4H6dHRrb5lzNo2Q46Dr/qy7HZWddKRtTL2zf
DsGohvaxDW4P5hJNzKyQ3GAlm94jOsv93BFo6PHG7UtwDtVdKdtAPAnNXzCRJ/8sEvFV1xy0UMhL
E+FNTqCyG2PgeauW0tccaK1s1g3/VdVKEGgoLoFBYGfiONG3OKJhh8rNIBYU33G+P9qItT2tVxkg
y907nb2/lbce9sMwThS8x0OGY51NqkRNi4iZzfpjpMMJWh4Dutu1kLMm5HDj2neDRrTQ0xvb2Rpa
/4QzdLShD0oce7bs+/v9b7+czWOfTtM8h9Kxj5tiQqY6jJVZhQ1S+uQVk/uMU8qgeWGRUGNxOB7X
6fGaHqGqH4bMMR85qcG1dgodeelQrUq/rO8m4UEQuJCb8yybanjMYu1ZkLmnRMjdL/iIRap3Pa3Q
o5fqTTEDcN+r2AmfpxTRgZicscdEkOlFgC6dRA+QedLr2mRR7aOfVZCfAJ3WniNHerXWFwJmLDIB
jsoDWMCrf88YQtdbgS6RPZhk6gWag0AHo0Q4q0tCBs7WHrdJlGSf4RNuUHtFWxH9TJQBU3Hl9kfT
UXpVLFWnHqOIT4S+aFGjj/xP9qVj67VTLsrIkDmXEst3px/H0AtDwS+y+/wuNaFIMsZC5mT0Nb9k
W022ky3IkFQfSa+mIEMaZ/XqqIfj7t56gUzggngmlj+vqM5Gs0Zlck7uyZeHN90nmvT4LO9QF/aj
5itWx7loPp14hjIi1zRZHojQ6KKSSUa5LES4bSxvBfTGSQuEEu9T+IO3BAopYqV1CFX9UxYEFbPP
HiBl/Ri2VRNQPoOx9X2Yi/BWZ9rkfvouDIm2S3CYrKZZNiOybLVSN+seQ784Ee/aoGGrR+Ucrs71
mtJVmHsd1HpBkZ3TLtUG6Es9iHWH4BM/NVv1nH6zS0212gMe7NyXBnNLnlcHAHK4PcOKrfupK6Hc
DGV96lCP5+lX1TBwdC63j8bWIognPc+pywsYFNU+laoWXT/72sKYioG89Fc8cB3SCNCbZUjoN6Pd
/u/hFVm2M5kVu3+aMPIMUw/RKs9b1c9/wnbtD743cVv91EfUTT7nnldqNgOuOlhdG/BK0OJ7GAME
CJtgg26ZdAsRKV06U8BY4x0AbQz61GSfFpHyWtlsjFyWXbnZGejNg+mz9EA2wV+nfywIWtZp6VzO
EjjAb2Q2ZjVnU9g5TZmQ5wUJY9dOyMccIbzeXAn7FVHhVldqknbnwMuoT8eKmGvXVdR6rWUQQF0T
2Ff9SnXrcCrm1fKmw9h4G25+3BNcfdHjW9MqCjCgtdd17XYBailPQg9zX9wcl069SwYsHTQBxK1f
6U/Fnkm3OtvjdDaZw5A7+Gs7ckee/MB0X3nLtvJu0IXN6gLwN7RcMpoukh2MQAv0aBkaLL0pZ/yv
9tJWDrAgyhszSzQAhvkcLQ3crLOdltfsH57ZuPrOs2rwKB+ikXSdPmtgQmcxHlXFKI5X+k9sJTNa
RSTW0oKJnWIx0CkZZmWjNqf66DCT9AAtF0hMH2v48YrauvIRh6T3QbRIrW0r8W4y+7xp5nmvqUDy
1ffEByDhG6Fq42uBP9odfO+5lZZp14OiAzk+m20AWfO2S3XdAbQeXFkXjKzIZDrL1YsHQErbrd6D
L4645RwQL/QabBGQlY4ELkWfGy65tzvauI9kgBM8fvcnc3FNZeq+Lv+zSu0mjy7+XMTBhQWzy+H1
mR+aDjHOU5IyEAsezWJlalOltCxcy5Tvdm8FbwytNW1mCu50BngZf73Ry0g/yMCeE7WKy3Ii9hTT
1Kv3DS+yTXhDLZFpWE79XV2xGZOqUHWlDAzU5SqnjAIicOiFbXZdcJiWlGNcNF0akD5SsfS3kL9i
RmAmgOulxEUblz327tJmIWxHaBJY0VX/NjNxwG1DpOZtTKRo+oK0HdCgTfkGDN+bszhOL7TsQFs8
sSDAIaOU0fmoA2w1FxPod3Lq71Q9MpEdbcUceFch1Xjmt1rtQ3gIEoeGFbCimJzg/w/QDbnjs5Kb
xSG3ShGzluflocpj02BQD8JpSdwkYfVfNTtXQr141dUbhNq801Aocs+Ik06SNMV7jiaX5fkPWP+/
YjYvF+hXtONI8XA2mn0oidypFYMaFo1a3dQbCkWR7G9m4UUjqV3N9WRlXxKVDF6WWJmf0hOUpVMS
I9tQgJGYiaj78eU81ii397Ec1pa40Gmkbn84JYdd8UjWB1AGosUWJ6EyXX8V7s1hZ4s1TSmWqLjU
rfu+i5eWRXPY9GhBaVjsuzf8mG3htjVV3uQ6k7Sc0AcywtX9N86IlFTxBx4PO4gObT/N7VkPW6To
4P7LuGfTn1KH4wE84jovz8GrDLmoUkWAPGm+ybCd6MMMtsW8lnub8L4u4B1sf5XnIJKZfeGdPLg9
2L+UP13ErnZYDRKMsnsVL0HaLzjaf7GeLwwSvm8Ct6guyO481PPj/ONUwYlqxK8VDvp/QXPfXBUu
dbF1xv8BDefgOITUSTZu719A0incg6Z1hYO7gu1acd+AFH/Ed4UNtg1ksfssj4iZxABkuJ9k5Jlu
+kztIAUKjwSsyHMcp5UlzW0Yvt5POQfiyx+rPlvW4r+N1xQYzNyHc744ffZAK+hCHHglJ5YbJjbf
jmUljQm33i0SQUsQ95xvhM6G4d+eTR2LW5guxF3PCFBfeZo0a+EZQ7QL2kSv8GBI0baFHlVPs+CG
Wcsk/oSsk7qvn0eEz6IULZbnTBDNxBpMTPKzOUEZ73N57+dDV7YT3EoeM+t9EUpQ+c0QdY1xKjG2
bq+gS5VtTiyy6W/V/Dey1Y6Prqv9km4QoNxRSiFP3wxkGRzW7yWOpf9XNBCaE8Z4s953T4zvEyPg
ghsJUcj+o4uOybTPsMonEOyO2QUlHnOG5XQdU0ft5vCkPh38RdEqVqLwPwiduVzKV2XjT+BfGQXf
mdRcOa+nm/+45Dur2Kul2b/xLvpqjSqDUSUe/XCIHxwKTPPWWOQ4+g95yH4bf3qUnvm+DuEASZRS
dwk3rnGxXNM4DJ8PrCn7VOxqGmvwO4t3eRCMw4wiuE0TWhwvDJPil85uKcYAkz0NRH+EbiEr4Z6B
SoAgu2+QINuiilsxL6EC21pF0IPFYVCHx21dtlA3iKh5UtQjocFNPCP1fTmuWgrapFh2yC96DBka
tat3RJ0CoIpCroQksJ1QSgCwAWp83xzlee6p3YcKlxc200ol3ILpz5n9vFINb0hwmPpxdZ4pfhRP
uckMjwmVdDhB1qpPEABH4VjjdlK1poAfXA1EqeyoVdtBPXs+9DN+fNq1im5Zsyaefbk4ipLFNR6Z
Rn9F3poZyrYaYtiUcmPkj2S++wKVah7rnYwBDug25XC+vSf0NWqIz8NN0XjZvb6GPtRxLCMMJQnB
MrBLu1fzBlHqytf/pcINi005jKPfxkNZUukEzMX7heuhaOlpqsrB2ocToxHkXyQXJLsqTnntlkZ2
6/E8EERwPbCRE9ObkBaHgTCrJnHMK14s75hslNoxpNKDlhxZZ/w5Ec389S4GR6e5nmCraP19TGao
/3cyYlAr5SeV4AwTu0Nsvao7EYcNuscM6hWyejsEbIKMjaZ3xp1uUZ5Um7/H5eZuQW3gB4/vOKRL
vvlKP40XxdK+Thewhh2+6f+Yd6XCRSHa01XDy1rTvJqinuo40IW5TcIwveLg6id6lXcgiaogXM6W
rwc44Pz/DuQ5yIFT/DvcjKFmauZ871jnBicP/PK6cQUu85sPrhptEPR7fzQ/KlPU97+Gmlm6VyCd
pBi8LIBi6TENfWsDDdE2lAvi/RaIGnAJj4PTP13Swnda3a6skgcR56lK5vD//GOn3rBY1nevhjl0
x20QhdqWFrms4KT+WSW4J12y4Q+1ZQLOPmEc8NPWgCsNhbDDK+bOy9OUKSEMAdm0oWSBHxfFVT31
6MHSLlXfH3h3/NfAYhfSqj0OUNJBUByree3Mrz/Uf5IoRhcBoD5VfckwrW8xCj6726ZCa9RLlXAE
YFcjUze0jvXGHEQkjIJDHNzM/cGFriKBjQbL+P9nH0rTGRpYY1u4UBDUwGIyOYmGultbdnpFL62a
VQGQfOZKiIokrJIx6lz3Kacm6UPgGozBVqZXkfSG0oS1HxzA264/nSvkf0I0WEkAf1P7GAjV+SFk
HB55Iajy6SCQB1oSBwnNoc+sUIIc9wEpQwcioXbEu/S18ueJkVkjbbXNYAWKWeDLvXtkUAxDgAKB
VKVzLB5rGfqW8lw6sHQiLgZY2nNjxVr9IRWtme7pOHl+gnVdb7U+uwmlbG0aNzKh2tdJd9yLxf37
zFOR5JJhYDPU5Sl7Gf0XahzV7psng4IFPcxaUEtPSmkQVC7xB4VU5ea1Zvkcjw+laFe201uTAjh0
NxrGWg3DnA+FF/qLul226b0ul3yjS2y9Y6KGkJFVX6eP06KsCF6d7Z4CZfdO/cYEBrPy1rJIO0mw
EaFtzu/VqR2RBCUltzVFHvJVpsvUFRQHkIZQqQlOk9XU2O92ITIoT8nbtVw04vnEYbCK5EfZQMSM
66k0tvkuYfGu95ytf7CkEJQt+tMSS3paV0nyx0XdCU2BLRLjgoAKjL+9be0kJtz6+bris3Ty0vXU
KKHY+hhikIAuDmMkIc3KjlsZPNcEwSupXGPPVrw18JE1j0nVlrmcbXB9zmaEws+IUpVRDCXtpHnQ
QrF8K8lm+dgLQUTDi1Ahg7H8FKg04kqBXhVn5LSZqOI/bp6VzxMcGSjz84qYqiHp7znpPKZx/f8b
4nSJTO/0rU3xX/CHTL9UiDXk6oMenn8qKwaB6ZHbzyhHeYKijngzeExRg1NInmrTplhcg3MbU3ZK
kkRZxaessDgJ0b5OLKRHddBJkqyfo8uePxElq7z87KRgy9y5b6W+ZcSChFByJfL0oJZcB38mTBJ0
PDnJONtooD9hal6f9UrEl1FelAjN720kptYPxmtKtKyrSnYZnMwvcAoMlbgFepKjCA3rOYV3iKqV
olrKMIw/vWvBcNMg3PvhqYzlthM3/eHiI2HhEzIUT95vJMj81GGaRUmk/3VaHdwctjX33oIbKZym
PFcejKO/rW+o1w5oRcsf7Zx3WEAkxkW9fyENpXbR5GFexd3NNDZ8LHnltzzmgBgyT1FhLUv40yaD
yTChe7xnyQgmj2JH/o33SQ/9HktaJuixzg7N5pHW8ehSNja1AyQUvnQYR5N6qoA7XTw0ScwkBvT5
P/PM+rXOgsr9NfFhDUPpDYAgIcPI2hn234FllelDwnMmAro0XHUf5r5efUdwn0Jm3ACBuofbHFv7
JPbyd8FmbBQWIkzha6WiYzfWmu0ClpgC65HaVN3jFtpROysC/bI7tLJI5dp5GCJ/DwRO77E0xKs8
nIdHlzv9ljYgXd1+2AThI6E/nnlTQ2uC1JYWMKLImFZiTsBSIW5wBvdiNLNyrrDm56Y6pWZWYKWk
SV4TkeZMrXoF059JpYwHXtiwflQejws2+1zk9rzIn3g8NupIDfv0YQGaFMKCyMLI6wvPRf0xOeg6
sn3boDfswfxZa6IqBj3hRk7qgZZqPx6QFzGNtYL8EZWt4WJDAbGbQkl78pWQq3Jf5sFemPKrP5D6
emv8YAH6kEvOd4MQKzRNc2/+JW+xI/QMJmSul6YeS4wmNNrLYK+1bBiKeLDRg1jnOiNyA4naFNwp
kPrWptJk3GClmU2Ot1MjWF5sflkJrcqb2IBSmaMFyFdJ7oAGiCFfeDW0lKBuLilxVsUUR+QjPsy0
hfj4H31wRLrsY19CMsoGvSoBPQb/k6cinaRDF7OSgDF5RhV8aTWJehLciYV07zNSK30GKE+KpHBx
zX8osVQod/zGmup3EShqMQytc3oMX94rBHki+mOfQdfjJxGuwMi3brkafIh4x4UGinFT/ukOSUel
c+UHcbpXdZ1m0wEa6sleBLX0bqWVNCnsAI2tNZgpSpkjX6UHIW+BFnyjSIOaZuqrPWr9YgyR8e2T
rE0YQFH1jMXR5w4TCiS/E1m8xuXV/fqmGjdLcBZy/sRoNaPMMqfgq/C6EM/wVldkr6UrBNF1x8q9
UGbg6vEBvu7g4QZuH/iu02stouO4mQJOeNbxiiPeSqv9dOJR0OkJO99Lpj66sHUx/IuBeZ2IvKKN
ePx8NxzLDt+Zih+Ah3JKsZUcREp+8qE0p2egH7+9tZGO1oq8DKiRDfK80GCwMySu4YJVMt25sdUG
JScxxYNCYWvdVzKbs6/ebZ9VI2RsRP7VaLipYPU7aDqMxScTZJMa9qA2wNOC3jcYe5xOe3RH2+t0
FtCuC+TFavjCY5nn/oPfXIW8sJ4U3rL2JJ0TytDMy1W+VoBxmW7XygrEIOy8ummGEF3kIlmULD16
a1o8hrJSfAaj/vYoPf4C59eiyUCrDAUzTehY3NzuzjOiGs2XtSZhOsDkRCkpWa7sOaDqHjMkHBAx
Uq4RsdQr+l0boKOujkrNp/i9LUElOFYLX1B02NXlSxGTn8p4/C6E7cXyWddjWRforOtGVVprwYMY
8tEuuEpMK/eLUJB1D4hQ1oQS5ph44zG+Kwd8wXoKCNDrOFsnbD0nlLVVi4IeHscPMLauyOdZUcXQ
6ST9Zc8m+zTnprJf0QIEah/vMieXpSQzT5lmGFolnsJg5y6sFHrBejEkkBJHHftsD9Pw+nYF7F3D
4PIQmj4KschEyhfVzmRoRFQsg/JjxlDGRv8qcQVad+JwhhZFbRKgkjjrLrUcYRwPtNe40A/wuroZ
06N5MW5D6rxmgI+Kc9ltkYyGMrDb+F0RAn9hmI35kpNIUUm1W+WMVEl4EkXQBSB6DmkVMjZiiCI7
+NIdO4gBKzln69smC7f3LsKoVC6IsLu+JYRo49oAIXxZopFUb4O+g6Hz0asAY3v05bsX453lliJC
SbbhhkJ1Zej4/2iPdGs1cLHGQBocU4j7QHGxjefHtYOmniibnMWM3Yy0GTciLXaGhmuh361Gx2Yb
8Zu1EbktdgOY4ApCmUFm8qougTob+Vm07SlSIaez0n/aYW1ndo27opAUHh1Al1D0Q/3VrD5iMVwe
F8SH67Lk7S206w1D/m0NRdr0eNf6qSNAhdz9Z5CHhwQtGw1JXX1SFJGyHPnpNbNxsyxoov0IKPFw
3dTAju+pA6WP6z3Ojrk1oA0273CKsXNkK2OaMdQeNNBgLt0q4rUe7aiHDFiX35BIrydEpusTcHKs
Se3s1McozTF+BnmUdSmc9NnXhv/O5zHQbD7fqTFDiXFQe6MokAwVrP3/MTIM3Bip3XWuqjVCUjAP
pZvZEwyi844GHU6QLHWWaQB84xYX6PO92mVLw/YG7am3lqI2izq4NfUhSxV2Viek9C4TtM0erSZR
SBT4MPeHkBQ//y/12d8MeJqyJ0qojPnArTc1dQCQGMwhJKvn4b8VKSRC+xLW5hCAmiFmMORcdjt4
LmRIYPeUS6v6cdG3x5rk7aACYD3wmrlPW3W9/cGDSefye5VQ5PnKscSu9Y6BJeRoYdHv3QBgl0DT
xldlBT6P+cX+QXIlEgxUotGjrYIDQjlupDutXUUzAVe4ya/Q5UdYgV7q6jswgL/TU+hf7QDdiVCq
vquns74NU8PY2cTDPDFatOxOf8pEKZ2MmGJ2m57JyJHXpyK/Zk2MErtLiE9ARra1PXfl5ieqoR3C
9nHz7U/ubWBoNlDslBGxAjGGo66DMwdSSn+wvp3wnpwrG46sNqWoTuYSIqjbMrUCs7u8IhU1je2i
Sy53xyX9EQNSVC1IT0AkSFREoMvhyg+UilFt3RqVTKD0wMQ/MpAlC3FEG2x2GidAeKhHf2sn9vns
EcUoLCE2rrSr2/bJ3jkNDF1eyMjaxFcKgHTzKQJa4lfswzvjSNdQXoGAywSS1gRI6zkHa1JYGtrd
k4cGhPu8kh13pZjjBOTzkZ+QGv+gvNNrUzyLmil3q1R1zJvtnDRjXp3xMvLjs7/28S2VTGqqCSUJ
3U7yihbEqxS806GnFDc6MTPhBY+u74MzrhninlPYoFg+TPX6L3KoXoK3zy/8eQLcEZde+GOuCplf
OwsCOSEJQ9x/kzI5vLop5v7aGJ+yurw0RyWWW7sBtAUfzeATdI6/2qjDzb+tgM/wffXmM9nvUgfk
uvRF8cEIJeD+jiycn5xZ0FX+9/IND1RzMBALCRtSsXRtkPTT9ev14m1aRuIaWrKK+y2SrEWgtyTy
Pd6KjUUKq7NOTu3LLy3/kizYOYAKq5O5N/vKtOAxnhN2rLK4AoSgYdXVeiz3JO9DWS1ypp7ZsY/L
QINtiWRkwQ4TojQqDfoIwjTs7LnBR85lFYO4WZrVGZbxnm1kFmXkI9WPhTb/QJpaA6XpOX5DyjzA
uYB76aXgJcI1rrTctoeGgcCwyPDFdOyOzWtyD8pACHKv5a1WL7j02t6ZTpD1BUnhQr1bHpJNOfBe
yHdlD3mClgOawrWVZ9mN5iyQ5108PYwIVKtc1XiDRBzOJfQOFOAiP6YqAZfrhGBzeHnWjYVeOeLq
wSQVg23oWF5/sNDT056juaIhPUAv2PB6skN0aYZCmZz3SewMXVKaPG0y5ulzv5QCYyNRaoSiTtgN
8MFU81OtSfa3nOCN5Vw76h9NfLr50raDENqb9hB+jiIqcvzojLJWdK1DaVUSHBkYh8CVtgipP3eB
CC+WXIGZhp6RUmlf9S45yHic/7YY9cw/THoRqrRsGLoOcE5RbFL0tN6sAKpxoxKVyjVzNecQEvh6
MbfYhDHh7092MYzMX7gH8650FXsAMCpYTWk1UoHgdP16cIigMxa7ZxVTSPWqgHgvv2/g+4kLXhmA
4V1MsgqfhPVHjJlbD/5SfhLyu3/zxKi62fGFD7kSLi5PxfUkPzR0Jb/BfVnT88/iFtaf+3mF9ngr
JYwFht3SsFFft83NEvOlitb+PkCLMk+ziZsb8qklJCRXugSck739ax2XhMKqyYQBtvxfrDCMqR2F
XUxxHFlT19s/LN/el8iiKH/3Pk6pfVL0KsEl07+cSd4dAwKWGThsnxu3yn2zWzL4rW6mMEcLDHc2
UYwDsQml6iQDJmGXcW9AsRR3U3/1h/H+qFyhfiQO/UnQjXTY31kio8pRGOXMPj9rVBhvjJ78mggA
iHCw0VFmJMWiubJOrwNrPKXpEdteRac7B1c1DcSNEa4dx7+NqkiO5xIBfFmKWP8AXkAKqOpn0UKd
hYNUS/O0GzdWcePeruLTo7liDD8JEOEplJPlOCuUlV0qXnznQbOhvw0YhuxkKSWT+YTWKEF3lg3t
hbAmWWHRtssJ3LjO9d3QHkTWB8qj+VDJoNlvVPq7BlpFxfHRe+UON2UmqUgqXQG8kbbNIxBjG4fe
qk43YVGHbVEsyrZVNE5iPOOGDI6x03bstytwrUXcgW0Qzh3GnFytf1adNhgWewhQXlA8oQGOsIUi
NTWuuRlPKSuW3GjvnHk8yOH2QoAvDv7AGli13taQ3XT7u2LLfJqFKv+rRYqaVYSO8ofJ0CvRVqfH
E3WYo353JgigAfogi28annCx58Uu0+ICXfEBfksfSMc7Lg9Q5Lb+pHVp1xB87DYjWUmViBlZa3Km
lI6WXm+4gIGeSV9RZ/zLEevJvVA7q5y/u33pucXwmiM9Fm+sbcZq/AAbDiyeG9ETS1Os6W7ciT3z
iq95HJ4dPHPSnhrnMD86pQRCoa1xCzaCi2SrxRnyKZlYBBQ2rP1xKcNDRIkKIAxWbKWu/X4Rfe3K
9WPFlotzcxfauQOfTDYa3MjdXZGwAWnRO4CNjNIRyxtNd9wT/kkNdd3OLosxMprHD50b+xJMsZrB
tmL2im58z2AFAxv5NFkvIrIi+DbV7P+rsuSPSD32v6NKd650N52iBOOxn0mp0VE+ip9kDQ7oWFg2
CK2Y6kJEAUzD+b832cyH4Qqnv5qlM8bw47447bSDp9DPz9g8IVXee/OsUolWhJggokYaPMeNbtNc
HVl9jE7OZKVU57pr7ruchdRBoPyPigdscKbNit37z2h9ECaBmXrl/ANpkgUdCQmZFzkdcIIbih95
/B93Po1LGEU2NSHP2zQqYyhaobT01jn1tuqyt59iHC9fKnddf0xlAefhVTzltKUJrcXEsHjM9TV3
M8MwE669tiD4D4+V/99ZdW4aphlvvXFRS9BqdPgfHZjNjxtbVNUJTuST9wk09J+saBo5LxQ5e2/V
xVJh0kxj6+leepQSPu3cU6Qw1TY2jYXtyTWRXEaoESKHEVw9iTn5anf8oA+TeRE4vJXQkDQNljGZ
TXNKbda/okDhZenQlap/oN2FCyLlIGWUDFun/v707IbufY0UFKBGUvjMVd0ttbnzsXhabSctZDUy
GZyZ9uslv6hRaZ5x/kxgBxaGW9QUdbWITsGQp5ZTfwhdzXA8jJJUh5W8u4Qa8AjUZa7RNmCzEZSh
SMMbIPUtXp3G4wn/RSfihAhEXYZG+C6kh12Ma1Wq3xtn4gZ0Rc/M2Wxsel+MQSFs0n6A7yLhltAT
Ed0YlHYYKchSA/c/FBYRBU4UOj2q9liZsjWhG5q2kISoZB75I+CMMxd2gUWzOgdcKPEwd70VCBuu
ucGxZ/SJVMa4S08kaHAIJdcqukI8OEcYsVJedtLtIZK8NitDL4uMqjqs9qyk
`protect end_protected
