`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hg4b9E1m5rWk/cX/h4qc89vkZWoPKCUKsRRttpTFr0VLu+w/IWoJBHPPBtu5B36GVcjkTZGomO12
FMgo8oKh+w==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Y8hPocn+aaaOWO8yr5oAfpokf9p87x/5fgIdIp9lLZwPvuY1KOW+mXria0SroxC2N7zIU3noGStd
EKf+2G6ixeLN1EYGY1xuLRFhGJF7dbeND0GTxgbf6jnkd7oSiqiaqdp7h/IFIjKaYHZjei0A3OkR
TM3+xPa3+KhNx4s5qJw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
vV2nVUHyZHNf7APigU0XuZuHYCXp6HRwl4Zp9wcTFBMtaqezFBQAxLnIB2TvNkSDrCxWru07h+ne
Vp+vbNMM5MGo8xjY6zwqzMy2FW6w+2sXHU7nTEI8TaspYoar3/fEBcmgXoT5s9nDN+kiM6ORWoJ/
4hISCCtya9bgFj1bC2kN6u24IDKRtjMT2V0PD4lOm8/dsbwdbvnRa+rYtLxbMzQdij5JWzaswlII
5XO4tyIenYFJjRpPPPWZuFko5Wa+XsaYcJO3iLJ84Ln/R0Xkouyw/IezfP+aM4WZJSFbvCyOtzL8
javUnieZ/BBWDz1clO40U2igM9z5QpauFXxFjw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
BeH8fGBLyXJpmuBrwVvCIRdGsKk9DQP7Gwsz+zB9yO5XBO4iRbGDZtLpNyO4/IIA1VVaK7RH+5rs
+G3Fl0xNXp5GEoGzVDCGNbkwAleZ9P/G9dpCC09fum+OnLpYTFKy+vuPG+Mjr3MIQhXtFdPlJzlE
BzJ/AAb9GcZ8lNIT1M0sRz+Qg/AenHmRsK7kd8h3JCGwticXnU5wq9kuX6zeOBVEaDHHRCBIZufg
Daz2Z+zqJvUSXBxGMx04Nmo5G4p/3BbYXtefU61rSZL/qmfvxY1INjAvI1x3lD7EZnEjhQaAQyKu
FFhOsCbHbXSjcjLYgxcK8BdZISOsx4eTHGx2VQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
AN5q5ufrMfguiDEBKO4AD1VrPRnR+isxsEW0YuO7cJzk2zo3Y91D1KIe2rZsiScQeEXiCKrxbiCf
PBXiF8D/4eh/KRG7QHXJ3GmqBFxAFrSXM2jss2oIDsQn3TomJRYJY8SRU2dOmKOQBfFdNZdwBC+q
BiFKvET2OqEYvA5Qr7B/ug/VxRgMiA48gNZZysCifwiHxvx+VI2khZgTC+Ee8XYwJ5gMWQaZbW9d
QjEmCFM8OTD3VhJ65nLteLW1aXdMVx/KNq871ywC5XXPERT9Qcb8HysvAdWLpgvujGvchIxegjS9
xMVnI3Nl8c8RoFpfI9QUy4LK+QySWBU7hiZ/Rg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
rbv0g7kDGmNEk5Ig0SwCuTxeofbEDVq9AzjFO6uoJsNvmaAl85lg7WrMY3eU8qpNQgPO1FrPYjDw
j7G9fiQlyX7amJ7uSeiyDtfQRPAPof4pYAD842BisUjW5gMqsQVoGh5ixu3Z3Gg+6xehwz+yVPzf
55XyJgi3SkhAHl5k98E=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ibqj0WHStKMG8Vr4J8lh/FKvOwbDQ5EIHcy5svXUscTGRzICfGeBVKDopFFfYVtZRb4wXDr5sKSM
IDS9TcWYAQnuJUOa6hX07qSPgvv1j/73+usSYomP2Yvfap0vSDF/oroGgRyOhvjnTfy2YJHKNF3s
ihcjCoxTv990HNkQKhVh43ZZ1XjbzazrLI1kiO2av6n0JUe/b9CynnSTyd5NlYBWGXIOb4jbywpn
2Q6YilGW4KGJa6i1IyQQ72whTF2dam6j+N17Dt/0Yp7hIf+iFjnRt2baLFwabJzrtnldpJIUnneg
XpxUNT3Jam76kcxEckRBRaIqcsnO15vICuC2CQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 334480)
`protect data_block
xBPknxurXEd00nyDk/iT6zLjE9NjQovI1dKyMEeProB1cJwEYWMlyCuOptdDHL5t+M6iPLI3yP1z
L7gGbZhinfJIVQPYEZVmRwO0z/f9UDPtGH7oFYOsRw75BE3+kUHGaPnHk6gQHXL6OZunxgxo+vF8
+dtVJwCikga2tJe7MraFiRIjXbBl7AJY0hK6Iy0wZEkce2tuz2DAc0L5vU2sSy2o3gz+RtgpebP5
uiI+gx5h9CWOU911fJtyhrj1DLpy/sbUj/EQF2ppQNWd/Ebma3lAAw9ttqF1+pOvItooxVqnMOb/
9+U+yQD3Q6P08ltGjagkU0+xES4wikeSC2ZsliHeNZqULWaad4GktqTwnbsjQHprFAH74wuaPEOU
G2RrXkaIRhk/e5khwiDOvpSwfHLSCGuRlYXmsl5Enzc254cyg0eCvdDjXqDyu/rVuUiI+TQhuzU9
Oju3dPP0cbhNCxZrTYLnSWE74XyVLZYSYMsLusCnqOKb8N74ddSVuXmok8ZIYlRs+eeNI4TMkMey
NkUsev263D0dSvoIHEJwzOErcT513fJe6IhHYmpHLt4ywgEns/MFS14F2fmAQRyh/xqD6mAwqE+Q
lxDVYAWRuCuS3eMgAHDOISx2f6bqm6Jdomn+/qgFuy5/3Cy2l/6JGK8CVssfQhlJBEE2MfdW5BNH
ncUkAvjNAshzvv5CO+3DeixrK9WbNPA6wqLLRFxhbGITfXyyalh4Gr/EbazjJtP28wOYIo5m3tZX
yUiKiOxIetxY/XM6Cz/Ob3RXn8RLSjZcwIMW27KLk2bgH+PVPnh02mm8wtNqfcTd0HVKrYqF9y2+
LB3iFmeWmPVYKjYgb8FVvxdJBXTseY+DohPavhnkDvXsnoWjR86cjKZ7rKQxCuOiTqNdYY5BVB1J
JJy3gNKXAyToOavX4OniSVyo7iFujp//aTJZ2vJZx1vZ3r55Xu6X5/3pY8FHObcBjNOyMWPRwffy
2F1i39/Wqv4eXC31p3TNYiiA5B97OozSlxMevtdaq2BN36FabFqkSLtIDfUbAKU5jMucRfny0MKE
7qSha4wAKEXkmVzJbU3nTkliXdUKkPyOVcIVSz+7yFwodXrO1Bzv12qTaP4e9iEUL+L1nZb2oNQ3
4HdHA8uWlV+lwgI0HhX9vC97q4xkjaDDyt6IHYvNhEhYMl7Ndu2ZNjrWPTbKfVteHZ+4dkzIDOOA
cbzmmylEQxCmH1LPt/htY+wAPfmqGzAxK9s0S6HPlDfAdv/v2EfBPNETGol+lWEgiEAYc0K5E0yx
Zn5bA+bciUl4M8vKeJZGL6hIaH5svjrvtlgtj6M1AAUVJGQzlMExM3KHlmQFdsWWUNK7edYh3rmX
U9aZ+OFJLCrQKwy2tlNj3/ZWv4AF2ziwbazGl+D3ggrRfMJcpGVtsDz3xOOptOHpyfyC1G794N/2
8gmSOs+NOH+J+Y/0eG1sSYUuWxlPxcV13bLXNao+fRB5idFJwoG7qQA5hjT2zmSb1Aq6aZgh00Sc
I6iUsQgv/u1lPcWOJOik22eFFnbKG7Dyuh5+6h1TgNOY/4RKc7/R8X2mG70QuOYawCyN4/cm6rGt
wUmFyYJNvKs5bjF9gySIKl7ahbY6txDOstLLashPCj7NlY/AXV5EieI3kt0IGMOG/NJyB4e7FXDY
XOtla2DbEOLiP6KqxhMUevA2NqGvc9LEggXPD1X6iki4Tu3Ma0rufs8p5RUg4/9fGjvYgtu3z3d+
CqvaIDZ4Y1DG9yyLzm/UGZS0D864slxv9lCZrK7ch0GdKKuolJ5qtwxp1Cl1W0t4uWmEUPOpgedX
ssXUOVTE+hEAcSzxz1FDLvT7rWaQlY2gXcCg9PSf/qYmh1pA1Fzw75D8z5JCddjzYHzit4f3AC8F
U1XuaNPm7qmC7FFUE3yXbkBcP3NdXEpW2S7YLbCjbmzCmdH3QXILCRAbohuPHq2rEHTJ6HKGBgno
PMBJc4HRq17cBEqIASbKTrrNzEhUIbaAzNpNTGwblifHGrs/+Lqc/zi0iMSW8KplwP1FbUmb5717
+AkT71LpPQhb8rmAPOb1SPIjkwDGZNQseWxIi/kWODCVAK255CylskayfFfJkmBzr6DZ6Ifd3MBO
1uJHBIVTD3s7S1+sF1ZUZ7QkY4/i/KbXidQbLOJVEGABWAn4DaMzBx8QCsS/cnmRSVFpzLEm7Vf7
uSDqhFfDfTEeADr6wVYWQGTHrZ+sFHW1tD2GSGbCZptX03fqvBZ+J20Fv55ByhtbgJCEARKkTBZo
RJZxdLjfBgOWX/tgjYPVYlR8FKc85h/ovAVTRxdZhckxoCXZQDq7qvOzpvrgVLbrp1aojyXeVQYX
6SGGjS6/GLEwrT8BfOsFhrvKg2qFXvnDzJFvg8tQhic0eeFZ+lEijZ+IrT9qOtVkLwtl4WHa0/VC
B5Cb2zhF0jcvLb2EX7arreTAYYxwKoNyic7cNt/j6Frar9B2uO18wa4EN+b0vK+Qk2YLwUsO6Tjn
oeBTL2ijkA4/Es1DhyAuKNSKDcTol9hgSyQrRRzJgJgdTT8FT8lUr+Ql5tvdAi/pJwypHy9wLlRI
VKsSv/XcZ3V0x+JIAkD8I/JysJcCdqnJgk0ZZDy77M1G/ZqzaojqWsw+EZ7uhbsm2XlKl0ef5KL1
+DB/DIpO8+VfUFHbj7m35cy0GXulO6bbDNYZj3mO0hC3corxvAy/CZEcnEBuz2qc9pJHTnx16wQ/
sQRAi6RxQm35v9ZlovpR3dEbdCja3COQYVXzhiFaJd6bjRHPN4U2cwhke/DxpzNG5+ClZpWS4KBd
ESIMOSWC5WIzjC6UJSxD+/4kytWpdTkOzo8iiQibZtsGHOjiz4TjmtFUTFFd5I/STo9jxuwJyvvW
s5WFPl3wZoCcKq4a125jAmL3gekhkyEJw7gjggRAxlOA5Ba0XByLKLcYQrnX0wO1S62gBULNSU+Q
xSMPWYP/lKamH96cALfal1b/4z1ynXo2bgRkuUPgD/V4TEErvvBJn1t7fWJHsHzhhM+jKedxSDX2
xdfHsTNH3QxREXcOsQSSA6jCM8YeQTu1gEQbPd6PvAdSmoHwJgBoeq71rnXc9gg9eS5yKkSXVmMb
1fcN3hBAE141+eRKBlKczFGOkZhuA2Cgn26bQfMepXHM7JNwH0lJUG2A0h+VQ5zg6MOcbb1pXyS2
bms8Yq26gqvybf3gYNjGLq/7aivTjryCHn+8rsI8wOkbDll6fWn5AeOAxO9mpc6XTsFMoo5hnbq3
7biTDTsWbOqjajSHdG9ilXtFcxZNjROxOnGVcTtqifx+2ShxF2+uqbqv/NySUqKpKoasAmazjxRE
aUIp79AKe+vds10QUOGgfTTnzQoTegcg2tjPf+GOtMyzno5YCIwvWzKO34ijA+iPkD5DllrKe9Bb
OHIc5sXrjdfbtrWPWpx2a73WxTQCoLjpHBSr+EQk5ikjiaDds0mvZSV9/EkAoDm5VuKvV5OWkc69
qgviZOYsjOyB5oKMgy4ZNW4WMfoQaF2GY3HXCmdv+/YSb9o21vHHh4Hii6uLMGdGJGhN4cT17wNU
fQXRfszY4PZeFh2yIE+ahy0GjCTbLWhDr/dWgzg2fEO568aZvq6HPfnqc07XAGfWpkPO9bsmBDCc
4LuUZNUkJ2DvwCjBJmjR2WuKSRUN5HRH95fD0Gx/aagGIhpe2FlNbyA6n/sEI2TKQxPjC1vhmOE6
fHYF83vKpj4Y1v8Z9bl1vM6blxUlVA2LGJEn6YudwokHg078g4Yc2NmS3jJQ8R71t0dgA1x9W6E0
mWfTKW/uaIHPPPLdspCpE0Uk0JHPayMX+8RosGheNQnvoSrqlQcxsYGnjuKudSZGHbnWbsz3+JV3
ogB9HkDQq2SxrvgxqfS7zw1uabPIvyycX6xBr9NuLcYKbC/yn8jeY1/pbQGFtNhZ0gBcSNGfu3MJ
x9HnZqPPx76JOK0xxHbV07mK6eDDdI9HHx/rJCifHmdSYoIvWK9tLPyxACR/M93FBStBr5yX20PY
xI7ibstjWiE/0SDakKVUuP2ZotOzYK3xo+xyh3Z8MsPX7HUQ4BIZb1Cjc987e43PUf7hWuf9whPq
DWI8UJ/evoToKJb5IkDBNcyIMHfs11CEIuP7PpaJLTfWd62s3kmFj/uDAFIg+Qli+mRDbTIwSvbh
9xNzN1OsRh1bztlUrtMUu5eBKugAmD/tpLvZEKJ+artcw+gdSWEquS8D9+lDgEcTMmntKUFAGjOb
OhdfEoOO8YCsDNd9j5pNB+VCBP2Mkjn3MRrVie0eg6lr1ZJ+ebxzFI9Ku637Li/9EJaFR7X6AuAp
+J+IYw2UnmioHVWoot03Ix+yEricEw0+CBdnyzkaorhyqRQzS9E5ZWbE1gHaGFvzDZMUuoEvjUSu
+Tb0DRaE+SWNmE54Ledwq7n9ELs2GnfiiEcTSqkmm6Uh+8LOYJDJzvuyFxh9lkS4EfJP2shjldKS
3FsmEYLOXKN/F6kLZgQVGVmwm4uoHwhhjqrjNjVZzyMez8iugCmBMGJfrPGRt/cX58btiyOyfWdR
1rido8QiK1lBLa5RbF4VgDDizI+BeqmmxVOpNccR1x9LumReIKVxULdyQxdageS/XDwddhprhOET
FOVzsG0eCnu+C64RIfMoQm1y6vOTc8uPmY099amrKBo3x5JbGAAYoIwDjJH+rPIUvShf1/bTuykB
bNf+qEiDZBqd3iyyfq2QDTyD3M32/oKjirXwNNQu+85VfBmzWnQQeV9F6KEBNqIuHVhBXmcTkLz6
xmERTmDCJk4Y7MCzncicFDmrGMC1jqGdGC59dIBsmVT4q7pXsNFR1fdPYhpeWxlRh3AUImPw5UDk
P+zeGmvYehqlTCPUI1cxlf37uHdJ7y1363qK9y2aFf7NuAOQFXfeh3ugln9VfL8cn+odUPNZLrP8
/FHpZgXRTmpQLSY2q5MWuc8Z5PumBLjptw3u/nXlMpzyozZAKcZ0HgoVNvt9omKAu4ou7G8UJ3dk
l/o0Yqlug4wh8hYLDW0fnyDz6L1kOIeuCBEYDUfpmh+FudKq3rAn9u0fYgEvWZn0bKDkJPI8go8C
y5F+MLA7f2t3Fc22JU4KoPQJuuDiB/TgEm/gpmS0+Kl9jqyPOYMuyUwn3I1v6I8LPMmvNgMezhAU
OMrTvHUhW4fBnD264Q4bCLUUIqgTKmK395CPPkdFZ1AtEEEdE8PHqzpxytDrdVSRwuCZtot+Myeu
DfDYoFzTDU0zUK2G/pWILu9chH1RzSwBPfMBmqFAgSFT9NXQx5As3EPaw/1tUcFx0ZvWZwmClC+u
jO6ldtY90SV8tLNlFEuC24kd8mxeL3rrekY8uPl0FYKNrDspV1wjtQdTLLyCpZJf2xBZXAzvO722
HUoqjuWyiUO6rAF4xiuN6bVWm6R0k1YL0Gb7zfqcrfTVr2FtVMsJvUjY8T68CquUfeLv+BAEy4qu
OjZ8tD0v3hDezJ+p94ixEBGNOv/47O52S14rgfWwPz4NnoUUEu2z5SOAd2AMkIkGriqe5e1/Ft5E
lms/DSG9HSXgcEtDhI8LEra5B/a6NOM89hLbXylPlvPShNDJ0QjW2YhdRtoWrvci30kHDgfE7FfJ
CPVkI3tmrdFYxj5Jv+RpPe1CD000qlV47ee15vZI820Sg1jfBugW0Mh0/Y7GCoEZkr8Pc8wJv2Kw
PAuwvJYyef3qBY0814K+qv3iW+Qsw56oGlUNTyEdimLPvMvyDcWSlRLaCYG2Ib9hWiOn4h3kbdWQ
k5LaRcmqF/b5zIdfG3Pt4/6P4yoJDAvmmg7w8YkWl0wr6dGK/HJKTTVsMA7Il4qn0ChlCfTD1CPv
+LEogxbaJehmncXJE4Mnug4RZk8iyL64huuoiFeribpuq6zCRqdlalsxmFWdJLGlJZs29XNR/n/O
+3jrIB12LHALOWnbNFc1mfHadubc0uwL+CXDa3NGy7GOW1tZ+rivV7KcKk1VmzIjqT4rcwWLmbec
ThkJa9rKiEtb2nVr4Lv4IKd1jfULEZRxsAKixxga4V/HUs5XzCqcE236HoPSY0PwgYdUSHY+DAp6
kprvnhY5qY0hkeVZ4qN9KRUOF0Ercd2fiW7cWd3HVmmpiYjL9WsintiInn2bt/ap1BhYikbT+ZI+
mcy/FujdFFXqw683Mg0/lXt8rSZUgMv2LbUt09srULRAX14iszf1+7XTSU8AAXZKmo+QJe8+c3k6
XIyDBnXVaoPeGsy2rHIGABOSfbN4zKpYyFebNrJbKfrVdth6kiuIIfz48sRy6b8yR5trNSCTL/ay
ApleSswPsek7v2NsZWu/vCd147I9IpGcvRniw56VCSepVQsfHFKk4ORHh+1HGS5IlQmGgIQULwHJ
xysiDwbrgfV5OBQHWq/zbaUs3rqZvzwgZP9M4+Ml5npjtgdDU2wRWQXRuFNu/xWDctQfPXiF1U0w
ER9YjZscb63D5KtB9tSF4XsdWmp81HRnHhO+jlUILkZrLQgpI3qjOXphDZfmx7waStAiugUGCroU
2OqieooKhCk6OcIr0hae+MbwbM7ZSysY2qTY+fOOMJYv6ijAHL9MMRNz98WbmnitMMLRM2PobkEe
EIYjBpuUXcmOsg1O4D/LA3jn69sx+7YM2263aF+e9MjnS4jI+9Hv8OZo57d2NmxfADSbDb3RFr5O
PepePzjfjMe+6Hiwz3qUZtbjceFLE0+IAzc9osV9dwq7E55hM8G4ej5TKGSJrHcmaNm//NB/+GrX
63+UZAT+wELEzjAQh09tpSSblY5alPVeMs1IYgxMMsGFfXcJLVE4K/tb1ww1+IPmS6Tmtyyqhse7
jvwXO+Ry/MUs3MxVxlul/OrynzAX4gAoY5jMD7SnLBfJQjDav80Kz6zBTjhczDGj457cJWo5xSX9
2WWrOmO4SuDQJP3j/nx/LfcTklUU6E5D5cKMDyMAjRIBBM3IDk5AHJ8mv3lAXVr67JvP6+z4QTqz
OQ3ynfxEQZQMDz0Ta9O+iPDHynhjFf6opFMScdSuX7lCEmVe4KEkSscmeM/cXR4SrkUqQ63FGHV4
aznRD2uQc3bD2OkIsI6lYxOtASoLRh5taRYGh2l0eo7Mfx+RCl/h3yYxSkOnEThDIDKyXPUKDBkU
WJBpnR1pAFCbX/rSw/nKMyqlhRWY/sqIJculfDof2c03ZQ/+FsgHzRgXWRQ7k72E/Fr6tp6pe4xK
gF92sPVd75k6ZCeTflEgGjZ5ziE1cIJRYOF0Dk5Ev2Zqx6ax6/hq299/n0AiQs+NuQNhiZpnhTDH
nimXO/DK7rCKDyKcNFKAWVbiDCkCAIUAPA51FZVfYMBpmwogn2YIY1bVD1OAdP1D91ZbzcGs0cbw
Pv4gADOXXhNH7cMCbbZOGTkhdRcusLV3GEWVtJy4SVVMKZlKRo5r0Uo88n+7PkhYqaAwf7hJvY4M
Hh7920vHUE/rL5LLAQyoyO5pM5PvuRi5I2cQjHZVLQA64tUKodw1Rpje0CTlAjg07FV/tyhG3EL3
B5tWRZWZygZaEnwnWmJhA6FwMFrSHFNwpP7gyAASBH9Q0ypemnfdEd55JhUTVfOhLd0mvBvVN4WV
68aSfeIuJ4mBr8Ceov7YtaDDneuvdEG6h5Hv7VFN+9njJB0H6PAqC65hEIVkQgIXpgAHuwQFvS4z
OjMvHKmzha3H+EymrAkTIG6d8r4LArnZdVWSo/Pv2gyoZlISS0xWFA5FckqFLRR8sWMqQu6qq6xS
/7EC0EgIyqU5+RrCj5PcZOPZ9VhS1VnOhJ+xHhFaBim211fUQMMfZC8aGpoaMbt718zVhM+IbTw7
OFzn6KGpAVO6QwpaWc2qmsVnG8iKbtdRw7DGf1oo/GlFQLTq3woiU6FsJfGZiQuHaBW/33ip3sFz
645zvvICdyqrC43h/VBQmcRlkCVwl7EoxhfnbvXOXxBAjXLDestPzbCkLgasJm7x+lfgGOsgWmWs
/mTvVx0al+rMi68eL4xl3CyiH81lyw9P6f1hRPqEE0GCF9NDKt7g3RLbmHsCbO2Ck5BMd1PxORZK
+T8+U+sYdN02M1B+cW+1sXPiZ9dVqeb1T30CTbNkRzrIsmulT3QKJgOQgRXT7dBXj2wudBWlLrEK
zk2oKZ9Z5+oYtLi1AJLQvVi2gFWXj5WeeMK8AQokDtQ+2Zfs3TFHehTD3P/jWcpPqEuTEiborYwy
ka9H3AAsoH8vlxksJpjKtbDMg3KzWCyBcL9KmQTKSXj/78VnNF0yLXw8sl/s3jCPcbvElfflambS
StQ7penJLX6rV8QB7xOZnXGBJd+oXjHqXZ4qPc+XiNFV3Lr2npowYO+OTSVsmmHekZryvQkY2WWR
WufQsXCiVQ8LarH1AfmYoZoIlzRTBzrhLFGfTvAZ6gvAbPV3+9nOSyAeODkBKg7QLcNIMgySVMVP
Dru34moKuQSzEAHwHxzRXQ3QTAl4ca+4rRqs61ks5x8CLWMb+pYrH6JB8KtBqyqKxQ9fcuRgAWUt
v4UERIsBciSiDHGUf6b+QePsdm3zenBy0wMvm16/OVXpm51MoO4dvc+u3vHgQ75qQdqfjrfGej43
uGMWt9fcWZ4FmkAuf1eJ3X8NqZDZUtMX0MmZpEUjd7iA5M9LQmhN9JqN3j2ODj6GZDW08odC0HPn
E4easzjy+bzR2oAASdYOXPGy9+wyR0WZ0IdP7ElA7F1zhJuUskTLMxxvUIC43gWW65A8ZhZvfG7l
vD/zEOcydpIKT2f0btNjkK7dK/lcb+3DRcRD4glY1iB8VAn0vxII5zxdPwh1pQjokXd/o7MNN9Wa
Qu4fy1r2+afZhUF4ayfcbINbJBPEFvkZpq9PSExIPNUSPlvErJKsiW7/3V5mEO11Wv0RuOhfWjlw
X7octXVfAnODAMF+rpY1So5nIdefdfEUdUriE9IiwmJGNv+un85pv24PCs1Tq0B/Kp/Qw0pQh4zY
01jRsU/Sv/qRtUgENHZimxPmjtVzeUxG7SQGa1ldkJPEeICzLNlTfStoQ3baG8qPxbITDP89hZFs
qPez/24qpXGtGJJJjc8PBs1CKfSqZoytqkTIujhHVGUaOjihoYhL+iVpnjOpzg95Qwo/CGEixbPQ
9phmbKBpEFN+PFtUxgVusGC8b1wNSiMMhtVfV0DqekTqbOx7JuizyX32qOfd6T7JLlmIG+clsCyQ
8vWpEHBxGMnz5L9EsoavhIFUglQYF9E+wJQcwHSRQwJlrYfm0YHXqVpw1YIFzCgSYRTrYA7didM7
7pIiLcbxGW9oJShb0n9dsBMjJrUxRfMgUPkdqhT7fCa9PcJ9ymt4+nuEBUjqswjHJUXVipEwHHgf
DcaFbrqzltOc+mn3Lbkd5o6PFRCavIODhjMStrYYX0X2V0DF5DCd+e0++Xt+JQFo1p4umEt/mdit
DtSRb5smWNZaucd+u2mS8w4iIAJkVYdtLzGSe8PmBfkYA3IiyJM/0GqRHBgk5/C8PjP/3ZBf5iJU
UyI6RWCafkaSEKd9eYDh4cgQsLhDtqaXHiobARTzAR7MABlbcY6KkhQTwKmYMOc404iDgG/01UmK
bpj92ZQwsddsGRihC9gWmmENUhVlpZ4lexRvliFO4NuYvxN0hqfp5z9PuMwmmwo0oaAmdfz8oXpu
B2Vhdf+298ZvO3Xs+Ewf7pGq76zwSYrjTMOfZPmGSSaHCzjtzKYudj2UvB0VgPG/4mIVwQc6Q4Z0
Lr1VYTL+S1tw7Hca2pks1VlRe6pmSJdjJObgOLT7NW5FH/OahR09H1x9YyjejP9AaeR0pURYFLPt
e07nNBcOiEJTjCGwHwn80sjeZRbYQ/2hPXgndw2uul+WPN+W6QCysfc85HgU4bz9BXuWpDV1gW3S
rnKIFa8ktmeueoI+boXkENuC609ufMHynSelmA2pPNYLpkB2A3cnB4/TSM0ZLOx2hraXQqr4kw+H
iYcRfnfheqk92jXusGgxfgVTFFo919gY6fcGPTLmvoY7mJZjWsXpoZS3gf+u/UuLwCXm/DNn3Xof
RWNoZiAvL6U+rUaqE6UJocf23AUocSBQ6UtnN/IVNq9+nzFcGpD1jqsqlkK7ZgC5WfmGNcO6B4kQ
pljN1DFenNms/f9RV30JOQQsua60SmJVmYAwJmJuN6A3ffxVIPvII+VB5Npo/s1raJdnm+HAvLmq
Ex1nTwSuUs8BHW1AujuZHSlPPVCZ6h0z0JsJUTJlZius046GH0UQNvOu1y1eX7bK03YxN7nILkkg
ZkLLzXeJMj5dobmOfl5A/2SfK1qvS28kVqd1bz5ruL39VeijsTRFyMDrA7EICHXUb0894b0Nelnd
3jnCWdVwqgIc8KNF41BNnF2YJBFjPN8x4JaToqE3nUg8XOwqGUSnre7bB6xZa7+oGuwIutsyeQXh
d5Dp+IcwXsGzneT8q5hjjh178JVrIGXY1TEwl6jx0B9flZ/3niHbjeNfJ2MWyxmZKjy2351XMrOO
D/2Z+uIHtVCK5nn81XN2EDJEtJflYBPHh3utaPjC2BalD0QjrUcpIULDfbnWxHgrBJZpJqA5j7iN
EAVWCj+c1pBk/5LC/Ae+iWxKqExP5klseBJYGA28SOrfxZN0J/HeQBE7327ZJL7Kk0P39fsDIDTM
5shy+s68VLVJs9x9+jM1stnEPfrHjAAnAvADGZUyTSaWk6Dr8zM1oC1W+0cLhL3MW3x0j5meLvGS
ltVj8micwtCLLqqBfv1Opem14A2El73Oh/pQoUKHWC+UBI49XvgxgAsVIfEYmnm4jeKyBNerQhd1
bYWGcPUdubjgRIq7I0a01eKDi4jxVXFdkK5YQ1tCJrEr3OLuVNyGL4YlNcGPwN7eQSGEIw+d792m
Gri6RH7N2nW36+hV0XwwJK15VxmKoexQnUz7WEGw1eAXdWa2XnQL7SMPC4U8c1V1RJF5ixuHkYMM
8XnJfZttdD4ybk4CnW732bThzT7uzjHwTZw6bkWjuCg3PhXp+pOc7wo4vnfAzqdWh2dq0V2ZEiEu
hBrIDR2dhxK8aY5P6eLDPjzAuTEDyyuzwyC+eKdGZKpIymLHXRypdjyuec4v6nLUQyklH1f2gKS1
3DxlVvoJXnbl5vwg6GvEABS+fl3LcuhaWeFNoOPmfYc+/NLl92QK3nrmvbesluLnLB2E0HsJkuY5
Mu2iKSP5toEcHnYWk73BYVerJ/r49ecaSYS7jjqzbgBxLiOjmHc256CzPsD/ZJSTeTcLsagVvCYK
M0RBqsfD34EFgzV27RRaSiw2qC9BMWqckYkbZqPq3Q+FQyy2/14vjTsszp2DDWVZPVdACg+/kjdB
ziXPfXn3FXn9KFjmF4ngsizXkx3TgfVNrpd/Q07pLmfvwyM8d3odHhVjZhSV+Z7+sRcplVKWEeC8
jxpgBDv+bYALC4r+M1KlMYA29TKk4shjReZRTbOi0C0WiwGlUXKazcQ4zk6wFaQrLnjpJsunZa4w
ZnK37OOwHu9GisK2enqA72+ulTYZbQ37089PjABQB9nyj9APMlDnLh0/6YCn1dwli+4lnSMVuVxI
9BkabKFocdhMZiU1li81FfT0BXd01s0+il7KFijijBJ/mafZE2YBExbn5/2WousgC2s76yiIHRkf
Ej59AHtzdI8USzHFezaySqPSBR0w0IdFfkzaF9nCDtBu9UeKlGHQ6XsKk7Q8ylPmLoNzRb91G4gw
+dYLLY31Ufpj/8QZpQtSFM56sExfjPY3xuSXrJlBEi1SSvkXPAKnnTVOh/oItnfMNvSUUxoO8xSc
oa4BUm3AW4Ez8v1mqwYfUwDZT9gxKeIiAyHXEk5Qy1gyB5WrlI+5YMl2WYKhmo2tTGUr5Vfg/C1F
CzFJo+2Ry7Ql1tlMPuM2bbfleCTwjUBJaxTSLL1KAszObaO4b1Rhtx+3mTvW8uyCLO5Kfigdkp5+
UmFLsfE+IibRPU2qo5o7CGlnMCXaTW6yGuF0fBh9SJhcSnpPKaaXchCVuLdqH8eiegErILQzam4T
NoMnLgLSRdswYDP+LxsVWLL6lp1blfj8hZEpAwxvO+04SuKC3p/wJ1yXkd2JcY+cDTJWT5ZkE5ik
fZuIYFj0EIEfct8zTsMpzjrFiIjiGSQcuIPP4OAgIUgU3DOjI35+Enh5hg94xXGPajg9/g7UPC7D
cmRsSz7vYeZ+DX8p+IjU2/qbcnpaTvfVhExveYiP00EmpBpixQVVd57M92hYBbri6FqaAa0sqrrD
yeCEY3dXbm3aE5rfu9nR1Qwa6wTIRNWg4qZodwo0mVY1efNoH0/gqh0V5fm82bW1+93YL9uFoKuT
87Xaurwzjso2Lc0tdVHnI5/fHhJTpWML55n+FT0PvtjrpWFcWdJRKt1W+9rGQypdDmeE1rGgqKUC
Pd0MPMlYc14VJRF5wg3Vl1s2xsn6X91pV1uVCaTeYHUO44Slafqss0lvakvs0dcL5G4W6rrCrKqR
23hhzd1MHfqpWHlgodiPyqDcP45UkkMKIUJWHCvE5sIJ7jHllOhQCpBDfqj4S3qA0OgI0y2LG/US
4H6kGsNoagwwpnQi+VKXTJVgD1DKGTEb4QWCHduUxqPyiIv5hutIURoPPUXdC2tsqebqixQx9ejI
9eUAWG+grBX0t6Fv1/B/9U92THU/FoP6Sf64XluZPoIMoPvLjtAOcS7Ktl94SPBz9JQx0uWAhTrk
PVgYBwywmdqBXpmTPZKxAm2fj0RYAeZ5RnVxiXkmtiMd6sezIci5sM+UDq0ENXJFuiyVccNLUg9L
CC61WdnXMZFVJnmkUZKZIUUgDuClt0NrZ8EtfwYHDcLZGvz6Uyh7JVWLcdmXxLNiPqTaoKjlvtT/
aAj5ugoTauqhOspWMycQ2ikzYzr/VM004cHZ1/hg1JtwYTTOBF5RRB12YipuZoDnEfQXrG2xFtDz
UJav1RgIFKwuPwmQSyEDWONSq4B2dgYPMKuGDk6vs6kC9S2eEQjXrLFTUsho6WziWEBYo5DjTFvm
8TWFJTid+GHcuj5/xtA5cCPBJLfYQSJ7AvvYeRlRfI5UkeUxQIbZ2IhZkRGM2glD9qTUrlL51i+x
F0GMb2hydO3HdewCKVxcYqvUFrjuIc7mtQT8RctNE5w87nQ7j3KGXK5BCqfJtAelRW2OLKZoVgaa
4usDPYRv6364s3AxDN2haZiJ32Za3Jy3TwXWAbWz1jzszt41bo3SaF4trIx0orahcSlQ8Ou3IC2D
NufoSTAcjyA8P5Sd2PUFBGQ9wHS2tRUPSs76MoZrDtNN7ug5BuLmhvnwz+K8xEjMgrCKcWi+4ywM
esSch5deMpdW2BdZuCmy7KCegEsTYahB02sZZhOBGbXDScld3aPYRqBv6ASkcChblS+D++P8K8Rz
UcVu/0MfS0jWqlmrVFIlg4/iq+fu0iSZ+O/JzBoGRqELoNhJ2Oe0EMHplLusc0gwcUjvbCL136eN
LQLQDRPXCY1LWQY/5LnoeHRA33yHRJEpFhBwf2EmPhzaf0/zASFwNC8RT2Vyk0HqFvkx0F39SL9F
dFbrs3djsrtFiTsvtdYuFZubtrFZXq6gz514f/X8dzCpHQy0YwNj9C8G/wWlfdmU1eGPeqpsBxGu
HPBH1116PlzS/n6z/cvrfstp9f0Ge+xUlL30jKKLgQ0cb5hHuo7vrwNl3Z6pqZMM/OvZTSwoWxsm
Mo8pdFyjZFifkDIIwMQF6urykzKnddLYR/2L2WZNI40rRCC+JCgP5WXkEypAoLoJxSu1DzVzt1PT
Yt6zeBfek+FWta4989RcX6Uu4eVIltsDJYRQpDobrpZC6/qEyqKCCSJzLX9nOJqzT7plLfX9C4uG
iRDIkUgawm9PMH0dcr9gGcnSfo1rRPSxcM9RlmEL3iUKFk5o1XvQBHCdaMAqi2q262H2dqQDeeNc
Iv4DFyuzvS2suchCvksdrEB7/DvcnNF8zxCOBE1g93GNXBMcuu1O5ObYLI0T/sTwT/ecPF26dVif
tJf6VRih1k/seGzVFPzjGnsvXrIxUzkzBtv2zklkQP//BS3oIJWLd7C5rncgD0cxbUxCJIHLG1E8
JBNXAd63wniB0yCliHOaqODuCesdZblMd96JxqYp3a46iOp6WhkC50ZNk8f52vnixGRGe8UoN4vz
qGjkaL//r/MBy3yd9zn4tgEGSboODbzS+Jtwi3zL8u+9MDlbRVhKLQWLuKVWauYl39IS9bl3M6ck
1dEP7E+wWs8tTYBUFfi8ZSMR688kE+trJ9v5RsN79462FF7YKpQEAhG9UOkhIacTYGAvXDf8QvjF
qhylymPOBejjrX0EurRlR6b0DECJhW4YZA9a0q5i6IHSSrWowzx9wc3lGD2PLKacF3tPZkMk5QlB
JUsdN2cM8eIFUY/ZXaPELh4iLp58g4sw7SKL9rshNPjD42/f8RnLYUJyyHsiKi9ztHGSYbkQdtB5
JoVmBKQRkXB5o/qzGWeUj8i+lp4UdxmZlBph2/JeAWnRNPrxf918CNMOixH50rBhEj01w9glhn0S
MXSuCpx0zojEra1YLAOr16+IN+sTG9Z10y8gsHst1oTMj8IA9CoyX4aXqSMkEraO+rW/axJ/Y095
MMiscMWtCDXmRDIEwoNQe0ORkav+G0YG5O0irPCkkxXLftuimtMTFbmGCJOdby3IQu8gESwGAXfn
YERq8lzpnR5G/s6xP2fBRWKK0jydudKe/W/b1QA34O8wKRKwWfKglb9ZrbD9/orCWrTKaJiFWRxE
zWYhw39UUhwH6HdquTLPUxHsI++BTo8Xz0D1lhvV26erWkklB6tRZs1OAhz37wuQO4gKJ9Usbnqb
PqNfF449WFS7z8XxbFxZUOyw6jwPPZGdT2ctBM3cl7FWZwDf/nJzAEes/O50CJCuO+NeIu35DKV+
k9pYhv9X/81X7A8zbi240kEuhieP7Y+tjZUihDK8xSXlFsaai0ugl1MURJvXJBCHKeGJWMojXX7L
3M9gRNXB42QnYOGVHqsUDpAK3/dEkoOwsFgW71/FD8FTLO6KlqacNKzAFwocAlLfzk93LHVGu8j3
aPfpkY1ulEQWZyO5VlHzVKkU0IXn3YfIKsKUPUJniVCO7AQwFTNS1k/OUG6zqCaymr1+cYtD5qY1
IK86vOhN4VL7Zsdl/o7pJZ5dI+d/bLVfrz9HBKzglRQwCNjXz8yp4KbHtEXVgD7QCfL4PHfnrl1M
u6zAvGWjoMCIPyMAJMYbD0b3I+HhAY8iPL1CXWf/BfTHfi75bhuQ6/HG7E32Lo4EhAqtrvc0N1FZ
y07wh8Qxq5nqi/oYZRuDSiAkWvHT97bGfZCGfQoGlBP54WGBtalF8e+I+8xDH2iCfPGDJh+NMMuJ
6AkqlUFDx9qS1ZnoY23e/9yii1E5vNdTodUtoQcSifyOAGBUmbKYkfjkcpVGfZvRo7S1sRMxSrxq
hLJ5PpLLtMsFkUNu4syXgMReAn/LsDoxGdxkSTTkqbEeiy93Tr9jMN7CKqDPaTlFFRU2YrqlqTV0
l3TW1c1vdDJiPkq9qjgYhjMV40eIprfvVW8HZi6emLCRziHcUayv93aOPwlkNOAfAj/dIwKOx/aU
OpRrgLLrkx+GZ40AwzlvnCydK5ew2ozJFTSeR2XeclwptK8Rc0S60zGvAS2ziJhFpyXXQ9cfxysO
zIwaZjs8/P22yfjGRLWgBvDKhLWRzH2Kd22Cn0iVpuHYLvQOpFtC5xKdI6kY21uKnNSQK3dWKA4U
91JH0a2xHJ4XQluL6Js6VqIVn/MPkIyHWBDT5d5fRycJdc9LLAJ2lgPQW+LX8oMgkZkZoJDrtTmd
FxyDZbCT1Qy0KJKd7DlRK0wGlgQOSR8vfZnkBkRR7GaJzlSjcWlmvlhVRGOn7hB/ll4hcjiLdmTo
qGmyESGPQ0PFyAVWfBbZsNT9TdVHKtr1HRjKawfCEsTd3MysDKq//p1s+iysCreJ9BBMQp7smBRj
8iDHTVsl6C2HVD/9p8UNYg99m/zt7g/CKg0VTcRDhfxQWDtCFWJbHVvGYX3FCaUY1qQSsptGEPJH
Ooe0qC7mYmF+AvPK6EupZ9jq1F1I0C+kCN1mQJMm4G2v67jt9q5yAT34uuTt5aCfFgJKRGmo5QmN
kHpECpeMnliVbp3GMVZzcMar81aah0IJEMpb/kg+MYxHuR6KHwcB/QmbJSuX74Ul9aMRA9ov6Rp4
ZKnJuscPhOy/MhjBqZqkGzwClDO+t6m/uMCWCN418AvxK9WRY0zkX6iHs1spwZpkIwaM5Q1Uws8s
SOU7XMGjzt+9xUCsxbdm872SRHlg+O2bjA2Bt8FfntmvUk+SLcSBuaHs9AwUrB4uvlOxmClymSZF
saSkoOeP5iu8hVPLGR+YMn7u9G5qmfHmnpX8TAfM1c4dRy/uuNPRImsV0Vmfo9SRn0orwiTJGO+B
KQC8IZeEikYY0tXdTGJFkAy4P5hQzNn1Jq5GAYslmAs+dFXjqmeusnrdmiegDFZCYz1uTBGMVXPO
DicSwfPdY2Z3uPeuxd/3TrqBx/EfEzD2HN2bDtqD5pW2hV5bO2fv8wyDk/Labg+rSassJwUoAzvw
XBPehsrQS0rjLKDIuFRw0ZIeifYfR7NHj7evDhqF/whGarOowhKAfxxP858oxtUqti09GlpJv5m1
gnU0SoaA2MfE2N1phMyEK8zE7FJ+Fvo7duhGT9fBwzsfd3nyNdPvifhVJTH0MzJQ7rgIN8iUaoxV
uR7pWQQlwi5qunFMrRmfAbvX/QEMX5Z92KE9gJm4m4Dz1mh7sf5SgHAagTlma8dzh+K3N28zpEEm
aCvARpTuGv2EEGJWpzx8sTHMt795HhtI2NQbOZRdHDrrPSXZGJHmQu8TaCk5PynJfhPmdhVLZs5T
COxuLJBeo8y6gkqaYm5eRTLsJ34b8gSSDeajF7wnSOnSMLtDk5uUSWeTnVdoDi0mEAzwSMQfoIBy
V4PrO8n99ki4JwPgIe2ozZoCOvsETYA49A2C1WHOaSyxmJueAiXkY1llCjLAvvS2ltpEjJ01MtYr
M5nKAhMRbydR4tBfuYxfwsBanY0nVGxajypThAmQojpCVPGjQebb7V+R2vodDNtz6rFDIUNoigwP
uS85cXb3LpFs12CKV04/0miK7dV86lnP0XLYhlCtD64MifL3rg3lk5nxnEkMudr9tV6CtCXLxE2K
FN7h2HzoViZsIlIsu7icaCtCD9QgCYQhU+NWdnPTuG5VMjRjoUdMYyrALS9VQv10tYsY/yb82uW0
oV8LVMFJ4phBFJzMwvdz6E7LXn3DdttzNgmxaCk6MXmTN4O/35ZG3sbHlKvr35jv3rjiheEzbX1J
9AcDtNsJZI8rjEzI5Q84dswxrrc0ZsDEPWuHAusE9jLBC0CFPlPAnequv0ZHmFevyM0btK0dMld2
QLdFJm5eOMc6VMtY9DeiI9Ej67rY+VVg5Oix8Jf6eEfGN5/k/fhpefYChmenc+Aiq5KD5sxAwLcz
RirNSM5lt+as9ZILA2aIieL8Ya8xibLD6F6c3xh33WdQzTKMtNJM4SNdgwqNVsIiowgqhEQCsx6Z
7fsCd4Y9tP9cs8Kud8jHqMQG7clpxEJokobOf52DzaovgcE+liWHAlMAu3p+wVRweJh0gnq7tb52
PwtgVFkSDDWIMmvoyTAuI0eGXMgzjCwycVQa4QZHtmPPQ/xLHvkjqluMrjGRlMIlK7EZRXulkbpk
aZEI7UK/qmYS+52sYvjfyGE9dK6RqO0MeaO6PptG8h//GDJL7czp4yQxnK1CUVO20ko56JNiJ5GV
efAiCrG0xnw2g563NvA3rWtFPMRogLSLgISC6zqBSBTzDVcxZ2hcgccbYZAUk+xuoxHOAO+Phg15
NGtdQgXQGCaAsqKvGVlxbk7IVwaKjM/rkMLKJRwxaJwx5FyQlm70qMenSn4P6nSjwf1GGXeFe8ZB
6ftKBdeFrXwDjNBp/cApxe+FSIS0WNQcFGmjqb17+NAsiICb/ajKmlgKXhIThkkG1y+c/kR8WPgT
J5G2pav02swSnCJ8nTdM6dJd/PHkTeiJrilqpGcNKG4wbsE+8rU5Tu8xNYzcOnWj3ZnNcRmkDWKs
bjTaWLhP/roJuHnHb3XWLB7MX7NiRc/+ZBMUtMCPcCikH6LM6VlIZX8v/iSbtdXcrbfdYbgis7UI
BDHvhckSqO8q8ENOrVh5txFtjs/BmK1g1lng5NSa1kfmmrFIbzX9c7Tk12EyAgKwr3bnVf9PL618
aZldOpWN0SL1dZ8XpOVQujUpv76QWFFEl+H6+Ck+dC8cVfUlNqohpsBq02XgOP97N5rrLkFa4A+0
VLH3RcpB5QaC2FHBOj85vT7QsRthunMNu4LDiOKcfhvkCelo0ndpYGIQbc9vPjSC09AD6j7E3wdA
PgLQw5TB4qsbwJ4/Bfmk5tsvtm+hsofDj0d71ASUeap6DWhwvU1TTQNbo5RsTNTdhuC+GA9ld2cm
5O2zkP6ASWOF+FnETY81FDz94tqpaWjogU04r/X1peoIVMW0bSM7SzqdFjiSj2bRRxpEmu8CVRkD
dLcBW8GutdIOxfoL7mub2at3XltraBefbRn2BmZHsEPx39Ewmzr07ktLUoByiAPlOlUA2CvkSpRs
sfl/jDXrPn/ihlm85F4l+BCy3mMHy+iRtrokaDjgbaCoeHxowFDDeW+SP51mqWRCOP1uvjqPECFH
Jqu/rgZdXouVPrv9bkQVZ6sVbda6BYxM+DuXGKqCf1JpQ7G6Q67x5O7aD6YK58Z43pVpVxt0AwUR
fyqccgp4rPVeNfVZEE9u8DcjIeVqtF3acV0+0Vb+Nu4e52ERKjw4O5BYupMwGJNYxeMOkF/zLlEK
d1+fvtx5erbGBZvNwjOsF0QRAsfaMMCkDbSmSznJNeeGVMVZ3q8TE7x06moAhHwnDcHFMZ1NqzpA
1Y40ZYdl6mQbiWMYoanYJK+eb2kWBXs2d+zaObZXbXS9jo2vOPmQdhT81kukC7UZf1b8YK/Zo9hA
eiglZ9OVmo07HnPQ4mayqyaD8Mj1YebdM4Iic7kCI400sTgp9MkgF12s8CiwBGgg74IJOMj0wJrt
zWO06I8vT6j5YRzV43klQ8QYjaWfxJ5sLxD849KfXbJG/PrzZaBFoYu2/NqIMG5w8hob//JuE3la
BbAZUNaHk3A+NBFNVid64d3TTLJym7nMi4GzkLmBVpLaJSEcA45MexI5+qdZssQzjdjs/OhwaqIq
mPEUnJO5P4pqGZeYN5HdGPyW5FrJ6cY2Qj7lrEIFd0tlen1QMBXCBLD3ymnzZTH1Glk0LD13irx1
uTNFRNOAKvPs0HtRMv4TLbavKezPZU3mzsgHl6cJS2YPv14x10StK5FMBzCKamZg5XdIpGmNbzzl
AOGOd4+A3Pr+WjvxFSyTjMdnX/thKR4ysu5H/k+JWgoLWhJoWLdGzFTLdB6gWXrAeW0PmfJpiASX
EN9PH00fQj06ovDQbhVnNzSq6yUmDXt7uJDWzNu8AwiNFJoZXB8gITPiXppPAbI8LJUZKvlV3mnv
fqpqhV4FBe8YJkZlPDBdibzlM6eG2XBH/Ie20YY2MlrwbXQKmjaZx87UkbKhXt4Fw9koxRtBZssn
DG110hD5Yn36ZEsrX1dvH/n5Qu/vcId3Sxa/zZ9FCGkNSDWtHi5khlxNxqwbBZF8G1v5RM4Yh/Lb
8g28WwK3/NObv9d2Q6wh0JesEkB3pX/nCW0oxVc/kQX+nyu701qFt1/BEhC+INyin79CdD5utzd1
s7HNdIafdCvCMhzTzvUxFK0VFvxLsGXFsRb4DPZlKrMOs/aAbus0RD2QE1XJa/dSpLRQ7p4QC9M5
7PyoGCjcX5v8c5Bh+3Og9QyZh/eJw7J282xe7ftXzp+o9K41cLALrwqNusc/C2Z2N8hEMrGsenWx
d+eWqnlHifUVdUzviGibS9o4FZZLcbsY3282O4Z/jkeSQ8Nt36jaGqtf8goTkNB8asCV6FN3fyAG
qbKlTmA6GwPFo/Nek8sF7iTokG3iNfa9t5GKdic/xmAD4i8Q//KA1uNydrtXYBB3NFwugeAWc5ny
D8W1PXEg/nzJJf8XwQ/DJv+rM3KyAyMd0zmr20XtL5Zbowekf8zh3ECX+NUAfAP/BYlU0P4yY0hv
MuFbCit5KDXGSMGCjI+reGEz7WJAVfLtQ71V+laSKk7yupjIdOjaPnMBVN7z7yLHgMPUZDS1Wynn
O74FLtSeI9rEuY6oI5mENa1/1gRQtdc3ieCmD2t61a2L8jsixKBF5zUd2Mf1e5TAHt5045DX4JRn
w36kpreDr5/qrdop1vtjjOUa67m5IwS52KOur6PUuc5BY96RzC9L7mU86ameEwMM8XDPkSpd2GRN
wZ71zrYfY/pUhbezMCZ3dcLEGnRNIR4RxHWO5NLTYwaWxBqOm5vcIigUeYFPEt2CYIYCQvAQdtyl
Qc+Zx6/rN1rWpOqgUVWvx1dDJtTo/3yYGIuWwz+LJw3MQcl14x9RCRV8y28jkoXfV7tHiZMCd6VZ
XkziMEwGBlv5Varsp4u8fF5vxWTaToE8F/ST4FA8Eo0tHmDlW8vS0Ay8p2eyakZhRFKJJ34GONhe
Zxiyztze2uhzFBsfO+1qAJmxIqBDxhkUnJVArnd9xbaSbWarLrGJY0exDK16PVQk5qmGKzO/ko+x
6xwniHe/263QYZ9GfpTyQrY7U4+4hk/V3OkO6Tths7qEB1GFPcnX22PTScUIxCJhg4nzdYHN3Obf
0TWQy/WzgrC7YQfF7D+k22PbjtfxEri35Bai1SOqNxg2pOIXiAgCjaFDagmCMXsYi153KkTCSnnK
Erj+dGPWaFQe4/AHsKcWDldCxrH2SC1FTS2FF+8JmMg+cqRgQ1ouTvZU1kGVFQIkBDNyLDI5mV2v
Wi8SnW/4jhK+Ai4+LTaIpxILK+jSrU8bLd+ge55bBTpLs3DA2du2feOJ5unt7KcIDUSrRMqm39R+
kuOc6ufuBDggbNpvKHjRyEqpOIlKmw5zwofAoamcNmvR8e49ZIFnzU3Z7luRuwBXMc8ThiuZ0zS7
OCQRHZBx4Lp3zwkYqJqewcdKkVf/8kGKwiRQkO7No8UUwWGpgVoL44OCZU1PzL5uluiYqYYQYAfQ
Opxg52zu53cQYEyLn9o1NnEH/a/YwTW5TVVjSxV40/BhZCAwwF4YEBJKX/tGK82zCNRKikxV+VrT
hj74323sETNlYC/h5UbgjSgtJ9190z9mC9mdX+T/XFQUGG2vFXuugkcEalSHl/l24YBv+0YczhV8
eKa2avK7DhX+xP3zt8JQixK0m/6LSQSh13FsmFnHd4hdCKklh0MvMeKvCxtO1DiL5ZfodMG8w3cV
6Z+cF0DmO9mlX0elwzh0hZ0L7QWVv4enRGJQH15WBzXfDdwb5DWF+PQVnmfgmWqQc+s9UDjqP4Mu
pdlXV6uJ1HpCPosI4jcDXvOy2svQWI1nwZRa2nfuVU2LCung+HWhI8C9/OEmsDDDv4VowpoWEMfF
uckyvtJ7K+wbF9omEnApCtL4Ebwtx+oONbpxXJ/li0DaKZ+iNfydEbjE4zxlYOIwRSlJ/RJd9KVB
KPOb+e8kAvRJCTRpMYZaTRnoEkjBIsEr6Sdp9r5bokGK812gWOlk/Ja7QaG/sU0L7OcZF7SjwWJC
ZKA6k+GYmb6C1azyRJUEFizMDk2Aa/t7g9ZRB8A17lJWsslRimDCBVUHP9EysFT1nqGwpMxoD9JT
0txNJXVnzo3LU9A+FNXBTJAwM4SqMZ7C8yKZyXrFqlZG0saKRwgahIvVRwUSqwrqk5H9v8MdlvCl
RVYCu7HJcwe7fllNCBjmeCWGF/hUce8oCExRuiMvpAoMJEAxbgMXe5lvGVXBHR97DeCrDaY1QrB1
Bbq7XusruXe2ViYIYTU5fIWAHlI85N+bkNESHw+u/ahfb45831KNx+Bu2xf2+klt7bIfF5d+stfo
gBaUVA9Jg0Gw1sXi0m7vDCTr8CFDfw+XG2NyKl3NyI6IPjRsBC8YT5LJ57ko3g2UOHt+DNebqdru
SWJ1NvYQVD93w5oyHQRrZN1QIqRNoDzvLxO89sgQz+lYT0Nlae0MVeBzJWDtN20qflaD6daXB11G
dVNDTe3l5oWFIJj7S0cY71B3TU+jlBI1CtynV5wmtzFIYy9A7oDSvl7cLk2Y5mAYENbtThFOF4Ef
47U62Zs2KkeNLkdcClAv+RxkM8ZCezF4ddJySHUGaZ3kwCvnA+cjf0Rm3U5Gwo4dCdg+TRfTKu+M
0pKKH1jBmLdr8AoQeUkZAdmYbR+WqrZ9xNdA21kHgIm2twQMg9nLiQtmL4a0MkkmlBnJZWvo5dm8
MtUnfedxOXdeZxyzPdNcNfBPqGbrxzsyIBriyjLAHCt7HQ1mERLLQLFuMHzPlJBoCNte0uiqEXaz
0hxfgynlP0Wgvm3uRahCqebrcPbdrIKfTQCBrs86toC34ak7kIZQ7orGXgBEmeurgSFaujPtDCPv
gCkOSNo2R6shAJgFXRDww2dP1OBdGIDXuS3Y9JZzdLZrGS6TEdbyOs2IuUISckSxRvU7RLt2HH90
g5DJ+wZLYWf55h1lTTkifuBXp/TJfYUDFAxCqiprYjxAyPVBrGRVOKDk5QH7ZxiLhzeD9hByu/ZQ
0LAB88XJR+yF83wkxmBfCIyZDE5D2BQovPQosolKJTBIJ+/6XV22QDpG88lvG0XiN9UdlzSZVdd0
6yBDuZ25ZlO8RsQ/Be1B/Nnn7fTR4+Oem9HPIWYhK8M00kqj9KF8nKLIN3bmOVCJwrebeKpIYqKL
Z4hP/OuY7padtNNgpz3DdKLnZMB9ZlY7Ka/mSZ9RNR7imP+l1JTsVTDvY7jIXIEE4qpMR1juPKqD
O/2nqNZ7RHwfFfvTvOm/q1T3RsEMCzvoiSFmjtaY/u2iWVxRNfUcdMF0xzY17aNzR7m4y98KCYsv
oj8j9KzBDu+kOd2yJrxfRZDbfm8ETz+lKVMyYH/ZCuayO1KEX/O9Q3ZqJt3PaO7WOoQ8LzlaYwdR
klwfS1WE4k8e1MA/B+FN/SMSk+COSGLDwIF7ZRtExs0abHkInXi9txAysAbHX3yyKrc+IH9BWWB6
l2bx7hsDXX07WE6LmPM+fTtthrwUmgFJY3RqZf79lmven959NaZzID7n7mblM51idmFrZxVbnl2r
LFV1qFvwFJQUD05w4OkYq7YybB9aRR8sUmNeRrf/LxYhdnhj6qYPPdeR8bORcYPnGm7e2xEDEPDP
6skAxTXQjsuYPoSRiJL5WUA3XmGky/NLB8WoNDq+4k9q1nIv5X4bcev3CP0r1tq0pievGT5zVicy
wB/Gs9zWO5sywQnoUyR2HN9cWPptF2OCfy0G9Q4h5iD9AFOd7scyRx9UzzuPXJbxqABaCmPn2TXg
/VphfoY8//FAqJ7Y4ctr5wMFSKujso2oRk11miltNv/oOeZlf6Zcw41mWJBAenhUNS3YLxQ5ysOE
g6orc3e+1drJdRbdGe4w+uO6r3wHtvy72j/qXAXqmLYjnrUqmuGG/VgBINYUHghZzaEKybM63atb
YZACngNytMbYLL5L8NjNHM5VQ+w2Ji1UOgdfYy3jW07RYXdQSVPFNp1wtxo6zCfL55Vs4i8M6F3e
MSQ+h6Mwau8I9mg70EYde2xVwZGXgJ/QTQ6o+qqhX8bzHPmQ2ewgbeRdeGxx/MmbDZj/o2JkXYw5
sIm5vOMjZJHLeuG2evqjPqHgc2VIFuoVeQKRnjIZAbTjbZstKA/2OB6c+JNbzRsncc6qSPUBnLl6
XCfLg39juq5BZR70T95lO7O4/svOnLEqv8X9C+JWUPnTOFhyKhuQzd4ltUgVzkWiNFWYKuM8X9o1
JxGN2JmlnNH+5TwslOFssMOTZ5uo2mVhOMLs/OmsTQujDJS4XMKN8WYlJcX7yhfesMfrzUhCPISd
v/n2t9h1TWOKY4T0OxgNdbTP3FXDLBNuOllq46/IPAg7UHk9fdYPgNeTqlLT+5y/wV4rF0aPOKMG
bpGF+zQCC1WFJxGeax7sqmjVwvMYxWo6U/hns9cnxQXsmfdXFg1CL63oDofOESXbrf8WUqFH5clK
bqjbwAnEaQ9G0VlMHqEQQBOA9ZfqZbdCpSCeian0/XPoZek8LZZTuFm5UsZKmJb3DGH7T+3/k1jL
7j22Ahb1/0/NaLYsLVWI4FX6QdAG6H2usiXSem9gNGtMF4KUBr1Ns2avSNjAg7QanZ4WYKNULJSZ
joW80/aw700XHRKFJAlwyN9eycy6JaAjvnKfrldf422k4agXF9oOSASLpJLwi/LfnyPOX+xNC6IA
5iLuKGuZ4V4BZ213+VdzcA2TbFA55jDqrSgbe5mlu4XWnoFlKV/6EIDHGkyzZ7hyEjd5Vtvz6PRz
mz6amF5yEaQAvNFjjK6wBqiE00oPaugaEM3FtJXN37tMrqQoi7NZlnLlGD0coSDLUXsstwIiAs2z
f5S4ZOqZ1dJ8gVXmCfSLDmUNgQt3hi1b2fAPkSSRFkcaU2P5hvpV1ukiWAkbGCAjeXeptxpp28pA
K5thAPE4wPh0o13k4/E5mpYjYdGf+uuJqFJorEyzc79mO6M/+LuyqndGdyepv+NLNajoKGxhoRxV
ejcmArhR13nwu3PxrKNTcZa2+uzLDABlP7KSflYYu3Ao6qXJXT/GQW3cfhJFrSEAUqUSmeazC+Z3
51vBRZZJp2ts+eAtmCiWEBstnE9CX9DD/CaR+AZ8xFGWnSU4vS+cdcP74XZ3mj8o/yJ1hmQoDHB/
4/qSVz4j82AtCVQdPXeH9q+H88uDGXdAZc8aHLzu2BaEDyBvcExnTMQt7uppGiLT4+aRc48Uaa4i
ya0QfCwMXrsTJDvQVsS2Gd0V6dqG8vrMdqWjgWOnPu6OfgthMbIO56no5lsmvhZLYVRF/gE4HB7o
TmnslmWY5qBLuv2pa9NzIRkjgDB1qbu1+Fd2s3S8/9E92hhOwy0PobnXTt8/bBBqsQ2Sur8/WFV2
HgCnTsLQx3dj+YOJwBgC5GtxNtU3aGXzDWZ5OIP69j22kjE6ktxgu7fKML1CapErMJyhbZTBXTBp
L+0sS2AEjWnzRrCWybcoSPF2zWi/jBNOV0HyD8MoMYEvyn9HsXNILGguvFZHbyQdhlF0WFals9gb
UdyKv2plfcPYQKRPj3HCsWfpQ3lzOcbODp0vBl57FftadFU+qfXH8llURN36GgSU3jEAT3+NLAu2
P4oncY4LsAAFhA7Zh+nu5/l94IA6HSzVhzUpEi5L1LFePUcxoXcux4ofK37bHjvIU8hnOezhv/Zf
YOmekFpZ/n1CWyjigVCN4DWyMnMNqB+ZAEos4l6T+g6xjEQBXi1dvgviGXHshFlMZAkVBfT6MCTv
mI27+1fJVmCkfJGkVuFX80kLyZfRESMBRE1hMfp705f9I16521mpAUQoJgqvXXJBExF7zzFtC5wP
R7JJQRaiu4lApbojI8G9bpy15PAzE2iZqOp+jIHG+bmqHZ8XH0WSVzc9DHmN1T1yY486vhD/AcBm
r/H/1cL3VQ8KURqTPPOVJibpYCi9EawnRxP+zDVswbGhvqTFWAiV/IsW066P+4lCcYN2UjeC02Go
MKb0ZTbokKQvyl4mBVOgkvAR8nC+rU2tLhtV6prYI00CgHvIEHgeFn1TJ1EaAzacLEaMG5y6+ek+
TH2CNTrDWDunWApxN8lKa60V1kus3GAbdt5EUThBUm3BpGX3olcZBzYrLUa1pqAaLmlrk0TxewwV
XLTFQZoCSr9PyaHcV/7KQKubSb+RzkMAf5rBNaT82OvRUZcZntApS+t3l5STBo++OCtwmRLs9qYn
uwRsbqh+vZtguN5/nm+GJbPdQzTcyjUjzK8TCA0BggiN7zEW+Jf5HGyTwWjng6TorFBTAvWFwpiU
r/ChE/mbLnIkbBktRkAfwQk+QXyechxUvGppuTm8g9Rw2zlVQwK5T12L9Z1dfhCZxKRFaCsD8GW2
fHKeSkNe9ksMEhOoMVv/NykqnJU/dLjxcyL/rnmTaLBJiFi9xU+uI/tkOeut87Jpg5hVl1FpWMUc
1WPhDUBa3PsnzbzQVnq0KotOPPJ5iBF4hCGYT5BLXX+qakIoKvCH+H8mhquRX5ApuKbjW9udnq/K
EZvhhLVVxczOayW3AJs67XExL6IhCJjQ2ZNHI1rOk5WtgK8+WlPuQWa5wF3lexlDZ1W9q7b8ECmx
XZgVLLwaimSWNlky0iuIGvGBXFO4TifyJ90KjzajiMTu99O3ApwPE79MaL3+gLgr5jYngAIZ8vno
JdRMI3HE8vgH8YzFjkc4S4inREAYmnIH2eS9fQeYQstYjoUGvS3WAhF8Cti87TlGYEx+1povDD5K
GaCpqy0s2zEjEYSqPr/klGSKFnH+vviG2mDPf+2mdXkTUyoNimwQ09a+l9h4X8cYiWuCSZkHabY0
b9u2ZLmZC2POjnzY1Q+4TGuTaJ9w62FUC5BhXFSOQSfcrMZN8tzFfFnZUoo+S8xxze7T+HlZ0t1t
CkR4/ub/BgjxG4OskDbJe7gmeZkYByvWBaUiG4GwqeC8DX8mBZwtnFeojkHUFk74pDJhluyCtA0C
tIql5HTHL30XKiRdBcb97+WK8MSQjrIRpmfLKAWlDmj2oa5WxsUpLOG/4z/ijCYFOsXxvqrJtxQm
zly18O9jTxr8UoEwWhPKpvSAD5JhuhGmboaCpg4a/rmgY+XXEVZhQZnTUgdRNdIKX3pMjgYdVITE
y6dtr8Y3h6rXTlgyYzvF1f8Cr4sqThZU/N30g8S1fIP106X6x1QPoIeIrwSZDeLBckg7lLCUCQht
9+UaXZRdhrytsVMGGd3uuwdg5xFIZc9f+VbhXqAeO/ntcGW/dfBQzaZ51MMCdeCI8/XYFC0XqaJq
gRXFnIcWpTfoG1zQYduHx86iMgakdaK3Tn01cMXSR3y6ulipzhWo3PHxIHB8yvQ/ekUR+mZfZB1L
US11hOW2zmP0UXRzvuM0/b+F87pIDOstTxcA2hJzRZPn8b3e9aI5qnyaT4GcGMaaKg6gbggo+D9i
RcMSMSbEsN+3yDN3MpD2jJi9kqo/4OKX+O50mrY1LhTDm5yDDShv0YBojrXDuVSfhWXmdyc7moCM
w4BCvND7ZCg1U74Fq+fe1AJRLT1uHJOl2t+X3RMabk/fEVcMZW1K4rBInnngUyhjj8Uz8IaaiMdE
4I8txx88/GfrG/w631hDdRu5JPjhHx8mWdcC7cUPHFNwYNFvOf0ie5b1M5yEbkBjNS0DviQa1PvR
i64sunqAgRJ9XH+dyFwAqCghQ43COj8AaaEzSWk0W2Pdlp+B/Btejy0E6w9g4jGjMG5R/eVaRYdY
WxsBAheP04u9v9VeziFsfoN1OQiwkr7AWPsYGfr2QroF3Vp5HbkPOGpzyJZvx9e3bktv7ZgEhnvQ
VrbUCFl1W3rW+HCqAMq01L0WVNFEoR1559hxLjHgCmS2GMCw6HspjgrChjPRMc5gBMBTbAT2WN44
wXYG0CVaGFpQ2wv5Ns8kmiWZkI6RHzEHAXcttrrwGNQuwN7BsZiHmNiPZng2ND3B44V+l9FF7cRk
78bKyzub9BcMIYxAcf5IEyR7BT1tT3pr/rQtOmqB4cyT9nh/x+RqkN0HgSU6HwayL5yekVnIt1KK
vms23vFFxf7UFKM4J8ZRmgmhrva9uKBiZw/jwZ3MSPoePfcDwOgaBqV3gJRF3xwOLSm5lqQm4cR9
+3ssmmwfTe5aVHkPYVtUDw8TRqHd/67vPAVdkP1WvxYF2PPA8RDzKfIKa0xtglgIV9Bv4EdPejw6
eUpkNKOzcDhGwrsbtCpmhBJEIPxMiyNt4TF2a20BkmyarGQSAdbNmy1PE27oBQWyCD95qldo3vcR
rN7YyKmN55Ho+eQ58qktWPjTLjgiDVPFnBkVsY7G/iCAFIvppXgfsl2dwr0oQG+lln+l9L4GVc1p
/v1jyksXoKksdkhafQTluDDZK9lVew2Xb7PMgQBQyc33I4hvZwpvgLU0XfOrNUs6IadslRNkMVhM
2nCRgkRnyvlnKMOjkqxSSL4w5yUkMHGqCAUFBEp/6FZBGoqnOkLYQiDFFVI5dHHYCTATM4icPiDn
87SrITZJhrjvVwObGypb2BMd0KQvX8mW9cVsnB0UBdCVeYThpkIGegA7Rmv0rRqjIKiQXRF8k5G7
bQ3guU8xeKJh9JQ7zcRUy0LaR98kM7I+DMLUvct7EzIYZijY/L8tCi4tOj1LB0RP5EW8gYiWDqzj
+1R8OuvLusCQLKOe84SBZSBTkY9nL7oYdPtWKzvLURVa+j4Qi36ffN+ICKj+ZDmBeM405mjfKqtG
ZURaHD7o26MPlqh/lsWbln/cDMP6poUqM8Qx6Ov2XodDmjIiUDr1QgjQQq6XEsbl4b1v+8E35hQy
OALAlLG776VeS3AzhQB0dZl2D3g9haZws66vMOAxdY6sJ66qUirMc+wkfcqRvqs5tiKpRL9FZBbX
UTIeCRhgBwZ3fr1AuV8s/pyg6H202E72pC0B403xy3pPrXZY/bpdlmLVp1ywufHa+RdoMeJgqCmr
0IcJxUrUdbqJaJED8e5+PwerBelXaJcyL0WQ066cxjSQCHRB9fTjWWhm2RZKaUl28BaFEaxFC53T
xkI9kjuYXGI/szPVz+5uSQAyVwhVWF1SfrDgrULT3J+u+TRrXP5oymW02djA3I9kODzehTOcmo+o
n/kXbGuV+WK1iQJ4Z1HGWp6oEDXMRx1wpao/AyGYa9BHk8Y5JLzoj/sWDhNfAqxrsybrIbKCtLct
lYoqly7L5dMn3lzxm+gLQaQByiuTcqeY4/YRaCz5ugNox4oKrAIvwMMktNXc3xQldusxaZKFOUK3
149C0h4kWT4UTNgx7yTsVqsOQlMSYMmYqvsITGTJJSlZ5BQWMwcHn+gzEzPq2y0ZRcZu0VlK0CYo
pqg+/wDYyumV7kF5otUSpupMIeOA99Fynp8OXZmFeVsWXUPQPv4y3oSVWb3hlPyUc9R03OTMEZqU
56YbJWcCJpnDY6VXMh7Yfw3UiFITqXN8tYfnnrUqLkqkl6r5l/3hIXTfIPH6nQS0E4FxRranq3W6
1cbl9iO4BGEN2ilfTMuyOPZ8f9bg7UZe85VPDiSBq+s+UEtpFsPjFDzFmgdEHOzMdi1MYUXHYleY
QeUp3fIuSOCCeDRd+Q8WPcrZmetgpFXmWxfgVcFGQt8qgr5XhMZ2+ojXNKnjs8U8+R/BA087sLE+
raf1N6OGlVxa1ZJG2Fv+BV+l4xEUs/zfCkYJzMHgEhtdRRUt1GZk0UVAa0C0Xj8GArarooPcKtSM
Cv2kPljSbPGObEVj6tGb6ypoN1Qh2w2x6EYi5yl9sosVSAdHSiOZcElrsx21o+8nA9rPbMvTifR3
mGV61XQedMCgO/+OWeZpH0E49TUTIyjqbXlTieVk+0OPQyNy4R+JS5AQg7X+fekMqjVtLsQYY3ia
yaITrC4q6vOeTyGTQQj9ZwLvSPn1sp+aWZqvN7fdG45DJKuqIfT4cRCkSnap9SGCGhcJfZMKjG3D
DzU+oUyIXyRY9c3ZYdVBPOR0t19gUDkcLaFL9nTvFZiiGPU4aiu/IxIJWxcFu/39O3TCPpfhk4Vu
beYgR1rmuJNZHt/bgE6plpo42g8qCcJiDla/JNeD1Rbz+97jfumByq+yNkIjml8ywcCUk15dEr6P
3N9g0dZfl99QXug5wvEN7XSa6KQpuPBO230tYrnrFEj3i9cKbpiKZjx9UMBZUA/PCPl0WlmJSEox
rj2W7JrgUTA8ar5dRCmUPksahZhe0uwXIoWJAGIUNZFgBN5rw3pQ+XtebMobcgj4QEP8hCF1t5R9
gasc7Dhv9+mpIVrXrXV4/fGoUdhJIU90xBGiNvfSI+CSyc3rn9J6vZE3l9nTNAaHXOaTplBON/KV
KUFxQzEh8anfYwpEv4jkiWFgAn/PJArAM6FgdtCtYEfC/lxDXctmHzRzylfW52SO+OSnifEPwSnN
4QTWGhipqdJ6pJBTd6yU/nT5T+wo5wrLRw6AgZFSVQmlXRNjsVMi+SUjPtAaCCl3Gd3RBXBGAsOP
09stj6ot/vIS04Jx+OVqnlUaC7LugOh5pTUgA56oIqjNFNglg7QZFjx6+HnnTN7weFUSZHnRSx9X
Xm3U/gUPCo/NxQFlCi9aUbGnN+9T9tvyEv4cnlj2cGfx3N+35Y+78l/r71PzRdTFr9ZtF6jIt7+r
ZAgTDJErZ53TqighZQj55VgWgvTlQpBZ75/3S9d3h7nB86jIJMcWCsIkkPytZ/oBozKbvDPd9Zcc
UJODiKP6Hlsu7PS9TNovN0b3UXop+pTGijzbPc6vxRoGKhrgiW6ejA44HEZ+gZb+hn5SW+hMcO53
PlJ8dgxdJjfSjEGRzWViYjuyByU5gStFY6Z8iMgu9UcDqh7AOFNH4CL9h3168HwTy+KmzQyiH2RQ
Ob9IygsI63PBBlAXxTh605ZVYhGnlVbuNlLFgDeWPaGpQMJDLYevdoKiIhRgg3wxwrHfAyEjZmt2
J7k3/HYjXeBfCaoSjjI85Rj3tb2ik0BiM4r6Db11zIRWCzHw+izn1vh5WUJzFL/YsMGkZc7kkdQi
DtxJhKO8Dsw4DQjfS/TXZFUa5kwt1JqDYrRRsLMZ23v9a9MCm6Af7PUBGxFLg3ODFADVeX9Bo6zS
K1BaqHBRTwxh+mzp0Lj3USE9q+/I6iFngpLOHVd74QWSlPGT52cKvfPfQH3m4Obaua1gk/S/hhyg
TrzsEo8pTL66hUIYwBM5H9xMWyIAbuC+aPjpBK94XOE9k5MlsIoUfspuCSVESFWKgr7dhZQ37dXK
1nRWj5yxQNfsZ0VNiHnHt+FWbx3hx7KkMeK37vOHVXWPOWBbzhbE36jigMTY6XTG7pbHqnG65UrX
g1ZHEVDx1ai9HNNvHlOVZZ+PVdGSdfvYePskUBnpn0A1+CCEleTegoGOgkOYR6j0vWnfEd9RyExz
D9qJM02njXqFOkGKrRV7PU7Nym9Dmi5xQxd8CUMvWvvUofzkZUhUCtl720Rom9FjmolRLkROkWHd
efUHomGRF5VG6xTfHNvYiodOlgKkAmmbE4UmKQdzfzrsA3jUL/ImTSuPpEtAoqCE8epskQVLy19T
LDQoHWEeavDnLbW8X3zYSirLU13+r+6VemS3bixXh0QJg2u4MTvP6K3g5unEEpDKlQuk7LAuw8Hz
ccOoXR9VPxMbtYTvzk8Tk4K6zEI/tWfnVodqMxD2XM5k9PCbfT7Ai4USqEpVgeQT4ZXxHioaPRin
Hp+Jb3Jxmk+7GXwK76LDciBtd2YBzebv1SaqxwQ1qLKKocpvNSM0bovtdI5qYsznmNSgm7dvhKS/
fSK8oe85QksmtglEJkFRdeepbOUno2tqjAq0ra1U3Civ4TM/+D6DlA419FP6LGlMIEFcWsXIYhkv
tWFpRnVdOKPiPRDNqsI2Pf+DY91o1pOYZkSF4dgITDcuf77PmF4aBhHaK2q+TEpUMQj+/u02ALfK
NdZOfJ52eB3muVU68Ijj0B/9YnWrBmWmAX8JgJNEuHly1fTQWQqI8k99FmkXNc12cnbB/EoH149t
eR2v3HWCRtwd9Bg1zqD4e6Q5z/3XKavOCx4fVyqAdcIfDn15RlY41DOBJhMjE+jxJE+ytwy+0Rwm
UP0s1ZPuNAheHpSGmVEzhQlODigEDjQruOAPLfDNYhPO+E9WBfUQM3bJguA5ozB7igwKH4cu2IzV
6saZRDTl31hHPMr4sZNeuavA+f+AnmYOzlZV/wncfZexyRyQW/rR8F39SUtwFhY8cOz5NgUuS/z+
lCfdcexN7u5GIdUECeLlejdq04Alk3guV8ktTsc8qI5tQ4Md/at1lYCqyq52oyaB6lP/XgfRzh1Q
DA23s3JRhQ3sxUUj4PutfamehPJ/l+9BjE2zwKfGXS5x8rG3GvCDo5LGZ8a2co/C6OWamRLUhNOW
nEI3wpLSh1y5pZdv30bxphWlPc37JiVLQWg6SRzoqgupKsQv0+daSIUiirRWxTYjB/iTZlSSKSet
4s+MSEc/4aUGiJEkWHGamMcObJJraAlKFGlfzbN5QJJ0iun17UP6An8uNgyRAoAXvn/RzVR1Z+1+
5ST+B2EVDZf6mkH9PImo3ltUduokO9DLyJqwQ6MnbLBXUm3RBFSioQOW0IsdzE5+fJ0/lpgOZPpS
lynEgonn0XSfLXEsA4ckQKbHbzq3DeujhxtWzkVzFsxy/DC2gfuVoraKizBuj0drcOXz22PkGFDf
jqIQqoyLi1wKmcvm/ePcECYZElqBBeJgb3j1PyuK7946Ovx/inPXwl1HATkQGSh+5bQ+ljJMHJwz
6XvC/vB0MR6TTLnRf3EQB9k+a10+syeXMMYQo5PvEV3Vgja8QOZO5FYwc01sV+0JAaBvERLVNnoA
SzCqRqhKy2n6CBM0figH3HR0vJlLNxGdsmlTmGc21xoZs0PlS/OkJ7bYQHh6bYnKwQtcO22+6JHW
SNcaGpcLsqMDPf5CcA+sdvMNgrwGh2jBV7AEToIcE94Lao3hDs6SIhDGoQeL9yxFcIJF0P4bAObR
Bqcstq0RtrefcQP+LcXMaurUC6JrulnCtTDXoH8qPNGasJ6RJZYiCTNz0unQe26F6+oB1APz7KYZ
+0nF6nfuPvh3DnxEz+nMudONPCeZ6jHzNIqJXbrW0J1+zbh5qIlvUfFHCmhLbFCLInKTOtJCQay9
V3Xk4hQcx5jx6qCuX1+uDZbmDACt/+wfAe7ZrDdoPIWqByd29Go3YR2kaaVwz7mGkYhhJoglGzZP
l+/BprtUnvVfWGeO3eCV5CDW9jR+uUZZgzds2BKHysKofVEYTOTeol3PfDvjWt7N07U7JcIcTg1O
DHgyKmzmL2Qy6rINacdLPNqpYX9/dlYGzvWtnZBvrk58iwdQRpGMj39e869FR+fzPAwWTgEUsjfL
+d9Df3Hjb3sRi2H7i9EPrB9Wba/7teAVvpUvObR2Q07Mg3JITX3/U0quJj9Pg4ljDXdh/6LfVy0Z
o4OSsQmXJUaCHqB5rK/fXgAjfDUo6EIuxhDKnu34057QE0igiddoNDmP14adI5s7JmdVsqkeNBR+
4J3c0Zuj+hHCfZQiviMlazfs5TO7OhHvjrc9+DAxMAbY9ePphTI5SvcynGFvss2Xl0R9yak/L/H+
EsDbH4wwbrpojy5ueR2jjsJCU42OXK7NPrWpJI9KfijAg4UPI8L9V8kJo80i18awqmambzmJkO/s
8ha8K1V0Tp1KZXGdll55VIoZBFetZ27yD1hzDq04KoXRReGtu5I29bL+8+DEU/r0aiUa8swBztby
q2Sg643TTM/yy1Ep4+wCtN0P2P6GjK5Q1rCfLcx5IPF9+QemrtWQUlFMUHbncINfbizUua1viwpX
4lqjeXFK7T1DkZmAe3MSD6QoinUWwboN38GPlLf1Wj/tNPerFihTAiDkBHkBkzlP5R6BaQXVmmiN
O3e1/AT7mpk5D55jOSCDY7dEGHlTBMCrQ+2NiKfzqB8SYlVYVafN0XkRYiHbbMHQ0DBx2SR2mCDx
m8dE2E2DChxT0g9uOojR3SnzLUrDIce41gA+t1vR3CWYwCqcqGLYK0jiqqAIBbpeUfd3ubioJT2W
lOO/atZBTJXXIta0at5e1S3mtb9Q6aEedpS+F9mr1KSj8qCQehcVmJkU7Fggz6Gv4YXI7j/O5Zjc
X3VYhR/ve/MB4BLSYAar35z3Ojsk4AlK99oyiN/Hae5HKfI9KPTqUdkf/d1eQTIQDl4wd/UBh5Po
ZhHhm+QaHzIHm5uKZraTzOBw3fxZ+V1VvkxoacNJCjAw/rmUmenU1B2jXuhGQbvFw31EHzennnVE
vwH1GYUtiaL0UWvgPgjJWrEInBmQ5Ef6k6RY2n++UdkV4LWRNNhWY1r3kjCphqjQYrmZHyM4rdQi
GREfJkBZ0AxykCl4ww+6gEKswJcyLAmVxOqm5grVOSqQSzJ2DsDX0DyEJIfBhW0PgODk9sX7w8zq
BAb/DdZAvNa7Vzi3l+R5h9pEGKAyMj6TVQnG/VVDJZdayu1vIUXN3atl8f9sWQRifw0pWJvEWfz1
lER9ETw6pVP/RePwFUV2MHgBQn87zy9y4FUtD5I0ccReWMU9CcUJV/7N2GPSZ8uPbrZfdZ4Iong8
ObdiQjHYgpwXyodM3U27KjxdfgAgnV0QeGl0MI7VCvLgMTbMNMb7OFfvrAxeWJ7uWx5Yfpn7ijuY
BDv5EeJTbuTD2/56ZRTSjlmMnK96UWF8OgiVo1ET5a4MV0gLKPvJdyZbX96JikQDPEchhaKIiGt7
gmjT+PpPp3HilmPiGCUu8hjN5HeCPk4oUTWz24DPjNwEEz/1IocAE8ddpdOqU8TVN3UgxrP0qGpc
Cc42eCOKuD7LAZESJGU1k0x72SAec47Z1FcIqEKHS1fJrqJzPx7ypvXJgo4kfY3RIpLLGhnjctYM
3b6jqgbSJu3GaAco2wTXVEBlEthXvctjhDbzdHKsVaGT/RjIMeTECD3v4dnxtr/7t8AEzMbbd4RO
KqVy7U3RPA7w3ruanzsaSNbe5ioLGg97PpQ5pTzakDtEL+EjE8Dm1gzNSRkP1PQ8Ocj9CE9u5irB
iXVGg/Mwbd1ooTANyRozwju28Qh/Od490IlbFziF/e9Z7WwyjT/jIoe8rHKU5P/1wotajEV29Vaw
KJb/I1vVpq2fvCZKnzbG5k0nONFuVctiFASbYRNYDiycA4bPpU4oKWaXondHIXaSOlr5DvBiD1xU
OqeHGeNfs9ps69Ber8/F66civmX6sb3o6fJ5zIQW3ywWfZIkSBEwEBVcUaSrmZYEBeSc/vayr3NL
PoNk/olUs2bSt9IIpWSWD937KHsv81WQmyUYcvamcDeFJs1XQCU+2sQyPqLgvaigaoybeAYhAiFr
U5hWjuk1S/sKtRsikYhuhCpVBJqiWhZl+wCkyokJJ1NcbWjIcP4HkzSgzlccfj5eLTzTflIKgi4S
j4B/zZRHiECUvgnQv8iCXGqLvE/faIGfmWAnnuWdyu9DTK6YLaflIjsei14qh5Tp/nxk33T9yA3t
aSK+59R4LhteXzK0yB+QBtsOLiNvE0rX22pm1vWv4KAqni/qIDzZYhEuzJkBSfiKXTlaacmNYsC0
JcTlyEbiU6C6bQeGkffFUcmTbQUb8TKloEYvlgLfjzFMPk7qer53EXGTYtXzHC1W5KHI31pidfcH
QRS8AC3V0AJSCeUG5gVd/i/Rj46wqhPtwJdtsBKIPudpOt3kReqEAiNvgvF2nkqdO3B2cRW7wT9i
9seauZ0e3P1iTKnsPKiMtlzLUtjKOkAfIET40rCKkfCci+RtURx/gitdeGerp1xSA6ChkVhXquos
xzHJdLYsW2qsux2DaWlMyR0gQIMMygiYyA77rSeNY52cT4g4fAgFVBTc/KoAiJBZoQhRDBwUIhJj
BpZagj3WECTH/vKqSWNY5EYjYxg2K3FG9ZgClkq3V3cuRQ/cHdRh8lyTsNqg6KDk/Qsgs5XofHtY
7/LH6CN+wEJmqv9H3HrtBiFFV8jeLYncrxeLNJ1kUsSunZysvG7pR7DNbcybdROjpZzTFyHh+65E
s86czvEX5mX6ouNRMjhKGNfLSNbzKRBlX/A+GQAN0zWXHf8w+wR01qFva04weOLax2y+cse2iLwZ
FbLGJDMfD6q49fMSTPcYWW/DKb9/YZsuNAslQvGwGajiZXv22YiQ0FdwHquFIHtyUDBvtyQtvOTp
Js7iQjOocrLFf0aq9IYJvCnEDcS6WM1iVtXJCZhLHeI4fLA3axVBZ14tsLMnvgR7LVL4Rv3nf99w
sDR2EbZ+JapYoQTu3TzkxEdJubwV0JKnMu2JkCsF+VrGl+E909f2vvKzHWu26oNbBCn8Rw3h9uAH
8j1FCENJrtVTm8NhW/owhH5S4vF78lE3scW5sbW90jO9yDpigg8d+T9AWmoWpQiQYIR7y1mzF8g7
fV/FghxKHi2V2MpbSoYfWXqvHXv+tlYABciq8Hx7oMDf1NOL06H5lZHZhYezGhM0ng3lk3hxYRMA
xHqy/HWlqFK+0nQ2dVERdkOQwoNRH1LMi+KtkyMyyljJzLajC6+h0TPubxyc1AUX6IWh85bw1IOm
JcSnnRZxUN+Hmi61vpnQlHrcnKpwYCk+iegdAnpkcYGynGUYcwMwl1tjNbLoW5v3yCIhEuqfEA8G
FGO1gr410S26Z+yfWwutU/FTyuChLRruKnqr4d1Vn2M8czBIXjS1+bZTVXmL/duYuJy6aeQkaU1r
V3mjHqIrrR1IcqoSQVJo6Ywb/giAtauTjQNvNOXgzxQbRfYazxe9VU04B6LC17wipz7Dv5Sm82iT
qhkXQAhy7IrC3EER8F11hEwyE5iW1vaofM9xBNAHAqCXnI1ofkY5lvLUj/fvLtNAIKjdW5uc2MKY
a2SMaVSq8bMSBnmz7ohtYCCnQtzkYRpFcZQHzT14MNiXPGg7gYnnupzCWeFWdEqKUvGzR6BAgAbr
iVoSB1bKUVkeGEOCruQxVnesrxD4y3clBkrAAsUE2BLAQIa0cZSsvAyY9aZCM5HNcsP7JVU0vKQe
LQ1/TaIi9KNsU2WGueCwuV2b15CwRGjdfR8cPeuP78wESj/BXsGhKGU3WnDOFiLuhTp6pQko8g0R
q13QOV2nGV4Zd1Ul3dH0Yt3xnmTp9q1ik6DpufLSw5f11mE/SDkeoSShFi0zKHJ9SgLo2J9UJeq1
mNdXxkOnw2H79jC3X5xo9/PakITYoHmh+HpSBo8RHIAcNFZ9z5d5FNcumXcpORiojOduUFDf+OfJ
7fnpFQhuMM/rNymc9COrPqPIFAos0lIsys04aFf+Niz9dAPivjIR9drWiDbABCGsRGPB84e89+ra
nDEzbnViXTf0MaRezoLFWyW4jBwTainXhcjVMEcL/fa8O6b73ZAwfst7F5xK1Hhe10KOd4byuabS
0sUzfxzhWXs/5qZisA5SGD6pt4HlyNlhz764/bBe/hVObkc+tAY//pQ4axvN5tluHu9Zs/viKSIy
q9k7x38lRQSk2UBNAd9ZIpfCP+dBrAE0GIGtNAF0uE+F0Kr6L3eM0LwBFBEumIm+0tV36KV8kfvI
2pj+32/vWflmF/5tvgHkmJk3My1sTDdCL8G5utCtnecs0T+TTs16ma/i1T50R8/oly3znBIv5+h3
WjH5zjOk8nXz0r1P4ETyfAGXw/669pPKV6bN+TFm7lydHidcvOo9f95RhfEnK9Yqsq+UxJcVY0ho
t/JfNy2Up0CSD2ORPy9cBUqSsrhvUn3XIajrvYf16Vs3XoQ+GF/DZpEmImwZ2waCNfmyUWB+7EfX
D6FJpgXoN7AleQ1dZbkI/qX/bazwVf8VO5i7hiFzCSziM5w+PP+RIAbwOl6xqT3VGMwmMzOVOiEq
Za0vJmKY/1VfsFiHg7atvQJoxl3ct96Lj8dmo20K8S9waHDXNnxquO6HPxtNw/ydT0+9pjJYyI7y
h4Gm2ohpaxWHhbFio2p8Vaxcb9PSOmaP15WTbmhG6ImqvcsL5pO+TqrYnQYBg9zgNvXg/hUunANp
vRlWCObbNVXgSuG+XtAipu9c2nQruU70J3ML7BZRgibPFuTuH4aaaHvhXF0ZvIdFPsdOSUHon6D0
TDiklBQS6mZX+avRbnG6A9ifu52Oj4qRPT6YO+jUiBcisPAA9edpS66fEMAd2Bq7j+RmGoyINWM9
bcMoNvEIbDo06BF6vlzwLPxYBpYbM9QDCr0zLwr9CcapCwcM9zV8Aa60QWjGkjQr8ALi/BCachts
nsI4LiAgN+xVdfiSPDG5lvcexl5uC7nXL93fb3Mru8S6OIkP/qLreDaFaFBUFSH8YncmfgHAXR3c
xEj3U0zLkYaBYTcrET0RPR0GdrXqaj71OBm1zik1RRboTmh392WwCfrKmvGPozpv9zwAqSfN9D4e
lJ9RTNlZ/B/D3spSXMyn4t9NjTrBnKqS01kQZBMYgJ6dn5WdkEdtH4B9GwwiWcwSkqEkUHmFE3lu
JB78bx44Y8aSsYA3jeeGc2Ls33SLQUDPC9eQe31QVbN2fp+ubEWmVFYWLwNEBqdrR+WC5KncQ2Iu
Yf2MUOj/K08Nc3VeAoK9HcjFrJZgfG4vxfPfHf8FwaRvXX4Tfk/ogv5yHov+v0XrZh6QZSnfq042
6rkaf/RdyK3E7bkVncH+RoVH4FEvxgQsCa7IH0O80iAaZ+NsxQAhzjWNP4ywzjSQVjv4+57gF72l
+MejY+BNLsk+Ux000elF1LIQlDT8MsRQ0qDvFbVL4dPoFjAbYDOIL8PLd50ZxOxm5FBq/i9o6L9S
d90FYYa/GYUeW2c5vNjlo1gpgRyYwzqdHUjrVDdjKQeNrUNZ0JsSpVtH/RTTZVTZgJdAGpFogcH5
tEkCbThdVe37S6UlJ/g/Yhx4SigAVMRwJfMKdbB93bnCbPUiVfBJ/zySyHmAkdL2DonX1cr/Ss4R
Kq3Zj9GexfQSszJfNTaPgKrhA7s0lpC6Nksd/g835idp+BU+OVhZHxz/ltW2SADy85czocLUamg0
KMAR7FkyVScrfQcPxv0e/m9unDD08j0k47yFJ8a1iMds9GZaGtnbrPQ78dl2Blah6p+ZoZvEjVZv
q0kGcqpBL1YxQRpg3veREjuYgWhdsKkQObQozJu9ggM1+0a5sbo1u7Gwc047eDWNo07lfpyeCD3s
xsCwVrsuLvM9rSQl47F3Prtz8DRuJH1HjS48dblLzVyEwzsZIC8dtUzdv59P+Hz9K3QaolazgGcx
jh4auA28v14a0heoO5yWyFN92XNoXdUxwkm9Ip4NmjCUp+0i8gxtWJ7Q/tR6+RchTnjCyAkt2EeV
hk0wNxHKyu96QX6tfa2QEk/Ig5Rus95b0W1y3cVVCqFJ8WaA19fzndpnmJDcjJVy8mehgQj6Y4Ur
GztqUO2hONRIfwXETb0ioza4QkCk1veC2xwPbI4BdcqKBagAe+bjfJdEJS3yXBz9M3IuEomhi37l
1IU77Vs7fU3/VVvMsCKSUPayMuVvPqkzLTdnk79e/OquYlW9MU3InAOg9ZuyrZ7kwpCR103C9eib
swJWUCuLI7AoZCIbKLyfs2Ojwhb5y61VrjB1HBO2Z1h5VjshDsWofBWV9hWSExMWN2foUyfE14gb
XRGwLj/RHevT5vFLv8n7bsLRpBSJeI4QT1Gy78wRrZ64yosCj2H+d79EMCKahLhJI0KTjGFreIUR
G2X//o6TB6OeR0YnREGYcFqOqHFW4aab+zCKCU3UehWiZZyYm5ku9tc72LUTfLYeGc3xYrgeMIVh
2pqb/MM78RXVUhteDzYKfAHo3QlrVlXsid6YI3qj4H9uehcGrkdun0CTIyWTlYr2w5kaGFDh9ft5
1c3f5iZJ8M2L57ETQoeekhHtZrfPfaHbmIiZgBOWHoHIJHpKafif1+wqofjrEg4X7AaZupsBodSj
PKpmXrp3yTLClberaV+xsKOGUQ+NRn9K4/KcNzoISOXcXSIbfsWGAQCZrVkJiTZ/rrpW8CjF7arR
Es71yPgWFW9vahXipQF8XYj0CbVqCtc1QIWhYHY3NQVvZgFJ1Gqv2bCMnNJXvxOFPtRHsPGwXQnh
+CQCLhpelZValxS+OrSGJ2hZn+7d1Ad0fhQe9IHpbaRWBeo+431aBnJloxjm/C+sAZHqe9kSIekO
bWO2sqtW3dCoH1a08uLQ2+kWUQ1fDEd/WXhw8yvsI/CbVhadzh9wPvpmfr3Z8Pb+VmD8OIPKLNhK
oKuL+hwhi0BxaKEOlJ+HmXAtP8BF1YO13ENt5PPuImAM49Woimk4SHU2CVNGmRd9XbfnFBrXcoCz
rrRkmN2+EoRRJiNtCD1WKcLkLBRDmYHLk0uAtISq/sNYSq5lvqRGyyNSK0Lk0tg7h37j4q4QrfHR
WzhVxtY3EHWejPvHZjXLJdJtneE/vVb7T2cXm0e9sBlrlq/tK1lcC+p6rTHdk6FtQDAiVHvVjUql
U98E4PTqXL8gQUBLvl6O3A5pL/2+eRvwmRrJbvumVrxJ3hwJ9yFyurC5e1b/jEtVZTOjhT6m/ydu
8uAXfdF/UddlGywq+aIdtselSsfZYiCUQo+NeussyNd7dd3wVlsSwLMKjlL7wPHibNGA4EAKouS7
X1kz0wdXMUuRAWGQ/O5Q8UfOOb3iEOulTSHryqJH+n+UKI1LA0bbVben830nbs5XPpVhPozD7qEH
+m8R6DuvbpDcwu062mqLcvm6gLULJ4ikDDh6pLEdtPlt4RisXlvJS+sUZ4yGxfRPwNTT/ZGCcbzP
Hdd1jB616dNePrUdF4FZP1/i94k8uPhZNevr2At7AfBTp6nha2Vdviz9q39FSPYC0bx+v+W+Rp/2
95x66CCuY1041BH+rKvzcb1K0jEkBhIwFSSNpxirPmzzMJmP+0qk5ECRQLoSAPl6JDz0Mvq71dTa
bUVWIKASSXbEWGObE/T2nsSWPUAmrWMzGo3c7dMzhAXhH/wQu4XKux7WQ67qEJc0Rl2gr1Izj8Oh
ttYce5ZLoe9sVh9GBcAGLm7h7XhEccWoDream+6L6W/xbyERmss7c6GZMHW1pKfCkl2OIoH4h2WQ
sca457ieHjzhMXGYQSijWi5knT8wt0mKu6aZx0OUFvaFie+Dy35VK/pavxXIu9lHNLfHM5nKHOpl
mH17hzj9ATAsxDD+dUWex/Ly3ZVGbLPodhIq5CLhmuybO6EFa0jQ7aZ48Tc/u942xvLkNVyOv8w9
cSz5j309UhCJdc4jLIZIBErVPgmB5xrJUDmHbcnHbMdjuxQpa99jH5S17/O2EJothTWRFqcIWLw0
Y1NNYpIHZ3Dd12S0gJhqcwqOHz80vUPku0O0UitVS6SRgZGNEfcD/82cbonacMxyl4SuoJogu0Hj
VhxwieESMbwm/jYrbfQjwm6nOQ0/RC65n+UC5/LWkeIdXXpaN+PJZjllr/5bcb1bdUOuAjknp/l0
HDZoEJVfk4AiL0idj8iepClrxqwAYtsjP/O9edwkTH12N3i29nmSJeJr8d0Qj13E9qSTTfCfW3V1
KP/3v4B7Vdenejdx1CGpCfC/TAGq+a90Wsiu65Z0KCwVFdRTft1dlpgRW7WNgQQg0Fdf6dpBzW8O
1hj1OHMg6IxTqBt/JTgX//f4omSA4uJxphjrgv34BPbghdWmrPkxgcy+oawQV4pgXC7zAv18iZhP
QmJpY3yMElDU33jPuyEC4HJ2Kt9A7Kl460sZRoOruc2A/Dvu3bzb0q2wKmPnFXGepgsZOW81X2/l
8iL0upRHIUx0jc2TFxxq87Dco11fod60UoJxsQGgXnhkEdyulhOmDVpeKNnaoTZClvs8Fj0NZrZK
YzkzadC3HFXIV9YmFJ/CwANpyHUKihb/OiXHEzayk9J3ucP6L0PWoGmxg1fSRt/lY2atUY456Hrb
BQ5DsWmm/41Xn8WFrIkhpfx4/A0Rp+q+wQBT/+xq6saTWxMVrywXQitw60LBQ7fZfdz3QEvbK7M3
h+m2GP7xts+tO5m02J9xmdfZ8OQlueKk8wRW+xVv2QsVb3DzJqZDicr9YpzdNrq+xFXwxtabknPe
AUXp7D+OuOAj7Fg+lYB7JmHxvmMzda78yn4LpXlI2xdOJMUAAeTJh0AGSz8TWCkbGIERuJZIG0tN
JoDsQAFZ3LDVeCdVLCXP2l1Bky7oDocmYs7qHXVFysXQMUZVEnMtSuBWpzcnJuI7j3MNFwXctZNn
dVAcsCY2bYA/pDGUgzM0dOjKr6ecdmE8DN9lrGD6HlAU9xhzuLAyfteM7zSHbg5XEshCHoHwE6hn
pe6ofh6IUD7QdDLHniTBLnq/GIEY5hXp03Eeb4Fx4ZY6Yw4bC55+XYuX4dfiUmoaEsn2UCzOIhnD
awYtvcltZeiyjF7CENvBnrD4dgy4YTky/Iic2tY1K24zxmPttnK5U28b4cMavIZSGBn0XOb80INh
kyR5myvJ3ltqlYluHkNt3jzbxLhqVWjzVRomzifIR9Sd+1NODYOPyzx/ofkhc56eo3v0tobRrxNQ
OQL9j4xFx8HDSKRb1cAV6bgOpUE/oPBN1wpuTU5b+PZIxT9P9Peh0OY781KcKu2zDU88Miyhu6RK
eo/TKH9GJbWHW/m2gZoARJbTMoLeUsoThGCs/hRYeQCsSlJJH/h/mBHsEyF8XygBkSY4HLtnvuVG
Ow+DrHfpxEgNSCe8NS3t+HkgWFOoFqfJXxHN6YI9oek9qd+tm1ofYi6k9HymMErhWrgjpeRjAwMW
ayD0tA0hMi9SZsed+gjciYC9GcNlMJ1fBxxw5YL2nn0GXbdd7z8nsQWHz7cXPfH2Yk1lBUet1uYo
TpGObB5sFmp9cpC4IcwSzsXUFJ9Dr18T8ffenWLOSSuIRlV+x/QaBtElvB2GlVy4dy7lJd3438UJ
X7/wvtS0pb9he0o3hF/BIginbHuHSMkDEljChB17XRtpW22eUH99cGjgbvH/1LokuHfRWnMHD8zd
cMIX1y3b0To7pxMl8HGG4VM2G8+5f3tQNi3bHPsj2VV1TCdxO41l2w0CErjbE/zlT+uXs9SqGS0P
X7HVgeU+66VZP1yjiyxb8L9leq0KMDykGPusw5EMnp/Ife0dfT/FYOv4nv4bbU3uEy50yWZL+Ja/
bAbDoQQWcNE8AcX6tby5ZXi/lqK0FpwVK7jJGANUmBD7qIVxn7tkoQBUs4tni/HjeFSJ7xkQ4QPB
FVFSgdXSO7Hve//fScViXM8exkJaS1+WwGWMOy6XljhU9jfjL92PA4qE5y/H7aQzrkYMbpmaNJoT
fuVjTajEd6i9Cqk5Aa3HADKAWHLkJza5f3iFCoXJjPfpiiTOA+1LP1dichhfWpjANZcgbnf0N786
A043pN+zcC0BXOQYhyljXgKXxPnv/XxRTK7cViGqX+6ciEV+j4ud9llGaSz8kxa7dp5zQCHY/Ef6
c4Mbknbz5DFtN3igz5eu5LXQUqUg0DqTm8Jqr74vbi/EA/OGlejtHDgtGE92/Ol4OfMyH5IhmgV5
ZcDG+W/+8qJfatQmBsD0iqhRaRHtBZ8IhgOE77uhXni6EJxYfct4/ZpMHcpn73yWdP3XYc0X9/+s
+z0SymtaEc0+ACHFDRyDPV9hSVIXmpHuxDcIPaVuY9BbSYPHHD7cUP4PI1Iian6G4WuhyW1xIrS/
hZK2UApLetvromrrHJWt+U0WyyLxTMMobpT43FjXmUbyMNxmpFc9yNYUPFwYD/OTYBbPvu41EJvN
Jr/dZcDAxybzE6uTJ7DTi0G8KGuu/JwOCuQHUAzb3H26Yi2amlYncjooB8yV5YBAtsQG2yvbfhnH
EsWGWtnHsL2/l84BcoyqjCTWwttQsV8gsRimgY1x21KsEVPIegIoG4xkHnSEXGpItNKhZfl2UrrH
Np1KD+c/WmV2znpZF0GSspT1+n4LVtZV8uWC9UO+hBXdJOLBSXw2X8nqLZuGI9ikQpurnNzjAlwz
09cLFFsPWxt7p7t7gdbeqziizCJwoYL5pLDwLqbmnQUwJ68qGmPAPrZ/VBipWgEbR/H8BAQUmtm3
NOkINjusk9dVBijd8JFWOZK4+lcg70zzqLl9R3vyVr/e8HenHzLF3Evcy32gKrSvTe5Nu2Jis3zx
6Mv5BA0CpQ2XuagmxkKBuaS1P0rppQgt14L7SODHRPXxeRQHMLm6jrjj+nTPaIsPEIlQPVj+pkCt
Z3XItwH2NfAtULliYg257nWgxOy8kZiMZnxintyHqogiECgjQZWlad7aceZAgtiWTRMAkA9rIqNC
OEu8wS0SaLZuPf50tCXOzcN17VeqLQ3bitF6/WQzHiosM1zogLqPl017Af4bTu4s2RLTio/2wAgT
YrIyQUWESQjzSfXHN8F0NIRtwU8LOH6EhpN4nPCp7Bux30gYpNXC0cz+sSqZvutix1jlAN9cru2E
jDM0k/w2d2xPmxHHgxUmjAOgctPMg4j9h8Zw/wN2JQ8R9nUFr/4+BQKWHbBoYs58PaWwufb9wMWk
cXFKaZrjl2wGLiT8iSsPKAoEIBq8VfaXTGLKwHcDbzcK/go2PT5IHLnSdPgpU8k4ccpmJbeXQaHb
UzhYhenLf4eK6b642cjRtw7djCUiS9D6c2G3f8WEaqgBWSiNQ41hbhLoqGd9gPiFl6TABWoOKPq4
pcjm8O9IgJcTsuIsULUOvKHDJZkOHz5V7dqTZQgLXkymRk3fSNoAXkB0PpOIdJLXWJH482dHSUPJ
kel/gNQk2gNdsYSsGmJ91T7ifymYZX3coip98OXJPVHkyQiUKLdHw/sX1CNBL7OgD+hZvaC6y6et
bVQQ+zzrxFyQRXVWXw24q4n4LJAO7jmIhHHWPn68q5I/5nmQskrQs9dxSQ2vedcAhmYFYgjJA1j7
jEQ2uTaenv4GkE5Ck36CeMzG3TTJ3dVBGODQhoKELwABywJqkWs8u0Lf4JsF7t2epnkBT6jGJy+j
qXE/xLtzSdYEBxy+k/V/g2oR6gbg7OgB6O5URZh2GakKrhHPMmHG0yBM1q+HkfBv01Udo/fq7e+N
o2ikC5WKpFVUk2CE79EigIKwLI4fyHm7U5Hn5hJY2ZNbZChZU4m+riiVuW4MPkXfwZ5NVEO3EpA3
4Gd6nlfi3IUNYIc6vhZZWWT9hsXTo0b+WktvhMH78o6YScUjJHINCcdO/ZnDv2fdCdujfwJeuB6k
zrO1qXfLwi8Jkv1g0g1VmL6MPRDh0fBLS8tpSmr03bKko5AqocfA84u+/D+yAsxZ1c1nqeVkRGQO
aTIlUCFsLfzVIDvFze8SPcXRunaR2XAZR7ueJ3hhQuNt//x7/JGmhtGhl7JxVFgMmImY29JQ85gs
P+9e5mZKe3weWw7POJf9ynNKC6kYZhQU6tPoREbbHqjh9szeQF1PZmrFGBi+TueWBRQ3hB3M43vJ
F+TKPN6/RhUJjiKLXf4hClgpRi8Z8X+Tiorw7mKSE94s+MIMGpANJQ7aDAqqGTewaxshECBmt0Xq
zrllXJ12ujOsrHI1V8BotYWljaU8aMjx0V+piTf7rzLAtLqwIX2uIXjUp3sQxVU1WjXiIbaUPJ16
B+5DQzTMoLYCwdSIjxeS/pRJ2GSL9tgivTRizLft7VNKdHu8GEBd9svumlG3ih5br/lrIS9gJ3oO
V902EaroeVYIcJ2mK2T4TUuwOhLGXAWGQpF5ZCDSqirlN87gS6X7o/E3hubUONSF78Ij6ZOnkSg2
OznT/OeGJSaV9LeQTACT+/jczlk2Rxur5IjlTT5iQWaV4YtGaaPDfmWXXHQR6LNRz2qPcl7zCuBE
W4xMCbAoToGZwJZV7HZJbrO/Fm2SkB5pGPDI+8eN8gcV+kqe4gEirS1p9xg03YzDaqPFhKeR+zU2
deYHxd6pDE94Lrmi60yAc7BIz4Zg9TAY+BYobCxKCSvatpr7xvn1aRkw8+9P4Zf2GJSxSmsb+xmS
jKDPsnIHgNJEyzAMh8EG0iflEVbJ2O2JKvOHcA4Qh1580pbc67oZ9fN4Uud9P5sBUfhjssRDIU2I
QweTq9CXpTMH0NZmDYy+ejBNviekhigeRUI68pXAZDlq7L9ZrVPNIfvIGGzkiHooVj2xJW4TuLlm
ScAvzLjkoXaFUUR31766guOxvORdxOQHle0HYAFb8aymKhJIH2upGHfbyySLDetsJ3XJCwE/jUaw
FqSvT5geb+i+lrtF5dGHpRP0ia5/RFESFa9oVOn7MNbA3KcKZeYB5tJ8ooPnA9izg8UxnxXm2Hmx
rfzZc90bQ8abKRutJD+iD3dLD3EIzhLYSv4mmGJZAdijKNrAtR2L0ctOzZSv4nBTGEia/gxlAfPo
uPnNcs0zJu+Vf4wdUARMYQ1BUeDr/lHHclCnIK3sExnKMhOTSlq/hvURwgLEBlOclML6mQkTkIo7
14+Im86msrk2KWiOuVW9QZaWYaHNNQhdrz4ZNnZEcO3rjrXDCxI+WxbjAiH50mwI4VrG+G8gctq7
BkEjtK2xAa1Zc5YiorSBBdWYFxo7ytqYHqjDuvzpSuIfKgoLC63VxhfkisADdlBYJzIe3fYfDUTp
HD7MmrmXIM8MlvBToDan3yOpopYb7pMcszZx+T7pZLiUozulr3pw30L4ggCI1kWtDdomaHNeKLsU
+GKKrDrsdAYanfS7jie+7OOukua0j2J5xmaVOHjK0l1U6hnL+YRpWTPzj/+1Q/nz7UixTmjiy4MN
ZySV+cWdcFcIQLx0ce5fzmIpsGgxipzytGNuoyESw1kPcaLCi2+2YI5zDtJ3W8MxMQCi5fZ3Nydt
A0WLR2vrbn74Q3KLEJUV+6LNA+3Fi01Z9gGHMauS9pNUAf6O0Y34wpqtvp5za7HdOUOZJJQ949HL
Zx0cQDPVoChVOMkYcyygDsEaXOpJy3jCIdbyOUkg4msNoBMPSlPvGUAGeUDDpvBDst3O1S51DYTH
78NfX7zD57jBNIeexicrSli+wvvxOmBqkkJ6Mpa7fBpC9uhKcm2ntqxrhdrL+O8WRwAnRH069F3v
pTVs644U0m4PEqtkAa3qHW24PJtgkt4rW1vGyF6fjK3bQKnhdff4e7RBVMXA32Oo3UKW1qfCQ7Gd
SbyJ9ph6oTd7EzU/fbBem5gJ+8W343QO0ZZ4Ljphx1mdu7zJLqTRbO7QGDfxn7UBm9Xln35JWG8l
4xtc9ymn4Y0N0pAG+dtsdPSDNoCI8klboXRhEeDlM6ra1gHNTlB3OVQS2rzYcdr5iv1hjjDJ2fSt
0F8WUdEpbDBXTWeTE1d2xhZKpo8gZEeyZDjXta/Tri1UxkWaQQkfYN+xDMLB2BZoA95brB8aEoAl
NlQ672Xkgqdl2G3xtqmp93uUPHksaQXza4t4AkhO2CxpPgNwPtWNdkM/S/xTTimKGnwrwdUpoo58
ZVOOvX4JplCpeJNqcGhvxN6NkUp+N1B1bPhwD6TkHq1zuKI73SNA9aL9WOqzvgEXTYOfbKtZTAZT
/Iq5B1isjFgO3PlSmabvlts0H3bRj68uxBHksCWwMkFh5gXfZ9sW345k/zhRO4dLskPt94W4SsMJ
fFrS9k7ao/UxbAcKDrmllSqcpePF6391F/M1pKlLLWdyqTjKJQaNpAtG8EnPwsv3MIgBvWcwBqiY
KcVZv/LByyosghuwuKJ2H7J7D8Y8eXl1E0xccSf3tTD8HL+4Fu3hCThBNV6tdOl3i0bETthRDXxR
ADaCN2+kj5ko0vbgthB188vdy1FZpChQNOYnhfvZVAZ6p7XQFNk87TZgYxdtb3TtRWrZE7OyBkfv
JQzuLwc89jt1yX01sK30XDgM4El13gTwiTwOuJGX9m3SOdRE7OruHwcwrH7lMd4yqZ5e6HaFv2jl
/KLL8TMMHQj0+BHomzu6DIQeCfiepVk1Y7ZlsPHkGSXPMo/SowBulcPYNomft4XfC1wwVqajC+u6
0NavQtDvOIcYMpPYSTMQn95ddJYAwR5C5rop9C2CKo0Wx+dlryu66DpdT9jT6CnIA8xTZJczMl9i
eWAHrF17kkbp9Rxl2pXcItgqVwBC56N8nr81OFLaly1obkJlnc610nOuFh1gXgxoXq2ZKu4QeHEf
pG4aEFTKusFTqYYJXRWapPH6UoRb4AM8VYm87DFQzhYdOTHKo4f9ekXetzHR9OwdhDqVxy9v6j/u
8qB9VQSk1FSZzmfe70kPhS9OVhB5hAY7L3XcrS8TsGFynlpJafzM1v0bttPYe5xy8awa3UqX2PEF
zsESf8SfifDBaydE+2JWeInva3Ta++9SRqjmbXCPqCw0igCCVnM2Vloa/Co/bih5NDB0nTtTOutX
r4kJLQ8aTzzyZa2Mw/9SrHUnjZSzxg0O9YL1ylsMXrF9MYRFCSu+CdzO2qNBY71RJZHYrh9D+KVi
P38eX6z4QtYYCEoL50C5yG7+UbTXFx8X5X3qgsiPuivq0wMPvIDgV1tHrRCH67B7JYGmoFKvX9tC
YgpuarMS7Men5p9N1GP/OfHeyCzHEh1UE/jSszM7bkV3l3l6jYZUpjHW/Yk2wLfmMcIHrojEfQBx
mH+gncMc4pNH2FcZWdc7fMLwJFDHkt5Kg7Aw289Cv+VLXrXqp7YjfQnMutjsPa94KNiUUfu8e9dG
i4CD0RlbST6I5jh0wrPqYtNKduwVBYQos0szoDa5kwIIDed7b5M+OO/d8HtcQnKTJBYaaAwksvMi
VvWNCng/Q9RhGinHXJCMF8/cy+U4adl3YFV2qXjtE18bcW3A/vy5/uLWlxhFAyRpzclrY/T8jQDg
+5Tk+KV/uCyexz5YU9hThElOeoW7B7b+9wNXkJd/kBouviMOOyH16lH8IyJ395T62r0aN7H9VLS5
AARf0aEl6kvjp8JNAym3sKSUZfyprG+DLORJWEUKjnNHNlpezuE/ABptIBTqU7cFSmhCPtM+f22P
fbvFiiyNhtVPAmnaQBEaquxq1UZzk/QuPNNhCTxycnc3t3h0lixTY6TMqlzbO+3RYXAD/wUSGa8s
WSG8FZ0jVvJaLbksN0c8nYP6zUhcGjKjrS7ZIGBSkjmy9Jj9RLY3keFZfJ3KaTliZWEk0ViXak+V
Yf5FMRVnB//pXBabx3m5zZdgXfHg/DxKeVabWSEDb/Zsk5FhCvCs8/yGPCXLwu1odywXv5t7ek8f
pSAYBWrLauI2aFGZXz6fvuRRZ+aBHyCbmNIAkSQGSiryfNgetkndVeVHcmlf1ZLmpVAeB4ss54n7
X6P4ObMcRwl0ToK0yg8lXAN5Slm0/frzEVOwMSUHzCdHJtdjoh8vxLc6BQ+j5pj0bniNRu6+wg2a
sX5CzDHj+vgxQgm5gXENXlmD8Hs4WKaNSsl+/IIwN9PViwSag92RXok4FJ3mRux+qwFINgp8ENr3
IMscUPXaS85M1bxP9+2fY+yj1uAUkpGRT3XVCyFh4+AgIZQK1RBWOR9JrfHj5RtmoFxYXH/HThMI
U85Oh9lktYqD2wOETgTtKnZCMjTVtauraz7Xej1MPPJHlKNsbg0zDUQ+sbL6LT0E/t7/T6h/TaFt
1R6q0rXG+d+ft+QyHsFcjW6QMlRTquT3javCbzDxvV5k49yN8U5K5JWSWn55zvwla/MojYAu1+vk
sFrGBM6NVOt6ZT7QxRiasNbaCKskvF0qF2xpqkSehfDO7CUqoPQKaT6y7kaDfeHoySZ0V8RZXor6
BQHI4eE84eLAJOios/bPrBrqwniBLuo60ctUwque4NbLhAf1L1/WQXmDGK5I3S64+oIImiBKr360
5aCphom0qPapT6t/vk19/fYpIgPKE2vhRN0c977j+x6gUWmrEQAd4DoUGg74BjtaetxXwh73TcFa
znu39NpaAa+af/HITmseeSNuUC5FRjBMlm55YtmtUnjr/uQp6HOL66oToXraORSQ11brVRttLAAQ
hYlMaBlcHXmSVC68jqDlzoXZmqPI9UjptpZ0bhJFkRd2E/GiTUij1Xyy/wlGzFAL2feigqAJiQTs
dA6eNb3LlsxXgZFuyimDSushvf/zltRIzRwZqy1xuloTQFvPx+CjPHpl0B6YYX2k8ijxKxhvIcPa
UrlitAtxO1R3AKue+aHPvhMUH5PMHPqNxZJ+FUCHJAQHJeI7dS1ThLRTQYnZgLTZ8h7I2SIbW8nF
UF+wF7B5b72bYYY8sRCyZe766rebqyb4l/t2L/d0vXzk6yHT8VAUAygHLpOMsYlqwZB6QfLj/mHa
/4DDpWdHN8ott1lV9m27NeZARrGXbqjxGzPpc1a6bchWhVe6zLplhQLq/yt1MP/EIzyLL9P55bru
8qsvPzmsFaFZW5MPrV0J1skyyDp1vV5oZUnf1U/cp8zDJZKG+3nTUPNfPJQ94RKIM9ZvAA1BBy7/
4JyphimfLyPdV4uxsn5r9FwLIftJ4Z2vpIvYw4m1KVy/dCss9OxobdrkWsZbbYeaj+4FX6idFbdo
InnHkm6S1hnfGc4xA3Zoooh2DiBPOpOH0rUhe0iUvzZc3P/i1O6vQ4h21xnOTFta8jvmHb/AcnMN
XFCX6huGweb2PYoigc/DCkIJFemGf3m9c95lMv5vBpq59pV5IZpdYJemazYM1sOVsmrIcNMVbS6n
xv47NB71IZUgGmVgCjqRZ39WCxoJEQH8BEymD8B7ySqhlyl4TB6fwq3YnDGYdDGl1J/km5WytD1r
P1At3H8D3JI9tRCs/Sxr4gAevCmEc5uE2DddIRuT00IpyYn4+FTDWq2SM7Ssxs819hcEd+E3ZIdk
/uRLm8nVVfPIfzsFYrdbvlYJYAwWboWMI0grAPobq6NkI38ObSTlUVfOzOeMqooGLR9HrRsYk7U/
AIvJM71zi2L45fiOL/aVYU5aYx5e/H0d6J1IJW26NoP7YYCi5aHuJAjkYgywg/WY1xY2lmODPS4h
X5l0RgcS6I/5FRmKFxHQpGeCvAh9BsK+hc13xbMvCcYj6/1Cn0nDzMV5xjghvZdAuwPg9NJAwlfu
gj6LB790/XgAtcvBaCmvWtBPMT14B2VWtSBK4yitPsYepHnzGja+e83R6C95gd3LxE3YEllV6oKz
UrIEI2aCpXGulJFf5ZyHac3w0jnRMy2jeT0+OEU79itIFhfR1dBJvYbNjV7IKsb0k2mlEP55odiE
xoXWPj6C3TL2BTy6Ch5DCOozhojRlkHNQmglF5EQldfeZNSKluc1iKms5tonTa8JoLqlkLmAZ5Jp
K24w8EmqsKyKBhiec5QHkpiTmP3nERtbPwLQpMebsuu63zimb+ConLo/TZHWqAq+LFoqd+K3u2iF
1PXkDLyfIhJJurzPIkR4g0o1Ru/h4XAkw8vM7kN6heDm29LlH3ZgWY9EVaQnZFBEcT8a2QYD3mQZ
mE2q+BHhABLjRdviPyRkDqDIsb9PE0c/5nOWCywREIpGWeZPMV3tpKWYGbYGTof3zVpRYN/1RzNu
Gtvk5RynXk2lqDChfyygNwt5kv3XFmbSko/jbOcHnCc7kgWkJd8bVLNKdbsEI+vDww7qYwI28EO+
WksKOtfG8DWhNVapTUoOCzJCG0t7icFcFRUFJ7SxQVtSyOBKUePJsgUzkWzTOTtA91pZdgidVrGO
jx3LI/qXX0bUvgzE79rw7HqS7gDs9PI6oBWQXWPAXt+2Bc0Pdu8MdBwADlbq5+ZjkHfeL/6uLI6f
GfGg4FB9Zm0GhQ9TRl6wBRxqfES3EJInD8DesGDknQDjM2ozFO0YNlYaORKN7PztJfPRS0989Yj8
QHfCc0FGo0w/3dN8NExrsglr40lF9/Yv0JyKUrKnQCmpj2Dy+qbZPj0FyhXpFn+1Gurq5Qls3PFP
JU6Y/LgSvnl9kY1OCtf20kQgqnD2Rn+9zlC7jDnQG30AVGWyGwcgj2uY0kl2f5pUSmKm+NMvEkM6
9UMT1rq9zN50Uc+omE9PohpVl12GVIVL8bBES8VKDB7gADnkvIrw3VEj0JdA/ATc8tlpy3acTurh
LuSAu37t5mujFuUfvBDYg5ZYvVjcrXCy6HA6C5RaM3KU89wf/BhKl9gTNKFwK2DqVZWFGfaGtV4/
ftm1/4hQY+SNDyYofr2PYxmO69WrBC1Xlt8YUUDEOlRLgg0dcQun/4Otrv3pIjVZUoM5QEyPqffp
dT6jyFPplmvA8+VuyFQzSCnBE6cFuGlq2bhaUBDBbWDJi6jzIrt9Ktr/WFyoZifLxj4dSTaVhQL/
qgT3+ealh/pWjeBEOEBVsNTdKz7H+j/urfr2YfsoqJ7ZIoa2DOHzDINRjtSj2HYfv8m5XmsyQllO
j5p9VF7eafn45J2R+LSYz9vUy/HT4se14gOKmz3E7knyFxjb9vJoBynnWmXH0vDdcz/KMtgdfHyc
0I2xUSJaZH4zcqXZ2LnBuO4TVXTwZKiyr8rwbFdIWNpHfRuWBuoD1jO3Jss8FcQbrpaTzPQihCNb
j3qnP56C4o8raCKn/MQBt8USLkJ9+elghWgNvfcThXaIe+Um436QD6En7vXVqzwfIZCPLmCleC12
N4DPpdGqY6QpFigGhg8EJUC/2Ms93aLAkqC1LvSPcSnZaC197/v2fsbz5In/Bf1uCnkx3Fr6B6S8
HtSwmmJjhPcZZLDULclk+iVCFWxmj7lLTM5R/lTpz9I5KC3AskYCo5tC2IRvT7ELPvEGMyNNFhjU
jhdu/YWTsef7IykwcrEDwTlDgfesx9sup+8CNbnGNdU6z3UmCrjPpF7y2Zfyi9R1fAYkgffq86Sm
qdqdU6bBOE0mcvKQN9wM5pEWBqzKmmUtS2EFkyf1repvfrahO9sGPJv5oNvdI3F4UzX98AN//7NA
XfeTfYcdcX8vXgWRuMRXPUYef46ZsNvLkUAzc6bMUDhD8PEp8am7GqJz+Hw7y52Yii0HtHwjJISX
Viv5jOv0O1LpT+UoUaOYJQ57oVmpWYHUfV5Fu+aXkrOu4ncWckd/LPJX5wogSAYAAkF4sp3Qjcv8
mlzEts2QQ45s+BKFri50KhFlA8XDwAlr9ZbSQyf9N5mkF9X4b7yvvm29vQx+BfY9WN0ECJ08VdSg
HVoMwoQ+80mArQ7FjYZXj3SPugqH6FepBpuMFDjYXs7ofhT32yJW4RU+8MBPFbJXFge7XOoOQ63o
ib+nkEsNg1WCjeTyO7Le7RF4bTH/j3UAXjinhyJwzc1xDihfDKugPYR5x92qQiy8R4QFsEkbcNjC
GlOZ/bYhjm9jLRC0WF2aGenXnr07c6AIrxFNVSMvcy265LRuAMiO41SoqTsudtKVG8CYyVWmR18z
UPy5H3rxbUiGDhlyLRSa/7oCYkZltKzf6FayDKsTC+2hSreN60Taw2SacPIo+Hr5LkpmJpQFjWWr
D9duwI9A8Zl0D9GmVyGU3SbirUdGp0JGr8dm5HlnqMX+Cnx7qlbfpMCe6600PPD8HI6IOyQTHZyp
EZeVq/v2TYxv5PJplYlsImyH1c32AwCqHGYvk2dWFYP0fZZEOrDeh2+vS0sKSC8GYM2MQ0826Ho4
R7pPtwQqP+0ysvhAumFub0DkJfEhWCces4JV3jm4k89CKOPOIa29lyt512FajSXC37/quaYsHLTn
oGW7qnBtgrQNXAfP9I9O6oFJZ2sqYGQCrtKTyu51Rz5dhKB5QRcUDQ+pH4N8QUIDmfDOLA4fuhPf
VeQMvBHu6g68Z8vgmTyM6fAZS3WLbty8N55IkPGj73W1KCgYJZeBbLPq3820a8VTWQ2F/JzkEBgI
39J1n1UpbJ8GNxegnitRMh+7Fz42Lzy+JvJ9zNShh5zK0KaFgLJpkjRxtVxgnN9rAZaiRFU06KpN
Exn06evXRm8k9NSly0bXe/am0CAWZ2zATXrU90ab2iOTozj2sADYTgchgZNCa7hAPoh3LFP8vJ//
IHwW7tZLZomeja0D9yrGucrG1wIck8rJ+An+NxGuPVSrcVAsPYGGsJqaLiQx58g/X/jdvx9YA90s
AEXKwLOKh2eBCw/UBt2J+7R8wtQTW/3CM9gzJo88TG0akznv34f20K6vSOCFmDMmZH0DK9PPjfcP
A4EyxnnXn7XkZq4R3DK7AKe7CYSX9lRYwVC7mbGyIt4yxULUx8y2SUS3KyhOY75FPuFp8AWP/6Gk
vstS8x77J+y6Ps5EQe1V527KkubYErbyEAt2opNzL5v6qIha0n7M3yI4aQDv0SAsS45Fzo0P9IlG
R52MVEaNF16RdXdxugIXaIozr1pERzsajPj/eUcYI2ddGnfIyoKV2huTy2kFNXlge+h1zv70OYQn
v6KW1/YWXxVzk00X9UPQrrj5Fkq1rMJQn6ZEs7RU+KKyw1ikxFmMoqBARamy7k2Pjzd6+sAAXjxp
EF/36xea40u7VWsTTp8147mbAnDB7h7H3eFz77wSdl2yQM9JAwKij5nBwrfcNEwLZXi8gd3QM61Y
FTjbUudgGWLE/zqYjcXK2eQZ2eYI9s64WG2L5ZuiL6N94XtD66Ic2k8mHRageeBoEBMsWJHgI23T
WR7qCzpPl6HomYqXW5bzf8qnU9iv/BOWDu9bnCM31z8WSA7oEzOonGpo9FetkfUdif0gwmiDhvFs
AcGmPPZqm4NTgc9jHxloDgbPqWCgQPkGfp9KomddKvOT19SnamZJpbHmWTRByArORi1vi0OfN2ay
JVnviViv8nvNuhQ2kHdIUm3xz+pkRVH7+SQr6UzlLlTL5kDvxWP5mxI7H4PLyK9tJD04H1pCMZci
67nuaszoIoNy2dz0f48hFNRKIPJqT0iaGcLDYV8AGdnxcynhg45D75fZ88yWHlDIpx0y1F6XpX6m
UyHmTgv7FKz0HVUgrhgnj5mPgkjI47sonf5h1Ifv/URVjvKMd15WRM0UQfaHmohRGTlVn2dTYkvF
Ffng9VTsIE0TaIPEdg+15HCA91hKYHXE6m29X7RhgQPjaZsN2RCLnEB3tJzxv/eULkJr0xCYpn+M
pxEewln5J/GTT1pZ/QuBCOuaKU+tdCfLV7tUaUOi2Lq78YMDN+MjRR3IXED4FBRnH7h31RbxrH63
cduPYejxY0bUwPufIJ5jSZxg1qcVUv8BcrA2whj0x2w9X5Np9WnxYPbioA5Ib7Z6iHXDqFNK0V9W
D5LNXiCJ6OL5OV53hK3Kb6TVbdhMT4D8Pxw2MsfiXE+tAE0qRKREXX3gYS/j60HUpWCdVe2VnKRb
6gj2rWKzDHW6Mg1MIwtUa6hWPHdi/AHD7CfhwRya52QIivoXnRAhK/M3z3serAyoORB665QOBfDM
/yXml+83srhyle3gmbBso74k0YBwxXws8OO9vFE59VbesJaONHu3fSb9bYEa+gaW7xnQu31p8du8
ZCd1UQ6JlGtPeuv9oAgM8cjOOQFom/xSURf4Zj0xyplH4HxMo62fYNt2tAXjQGIBzqOy1a4nFjDO
uT61RN0t99CfHks0smXUCG3aobCrnYvfshZfogOg2Mr9aEzTBthEQRe8MWEZ3h++YWndOTUqBULs
SUdt4Is6y/h4QLGaagf2F/fCb/HzVxPRbfjrx0+geMlbapJjj1xsrHaDQTz/oI3Y26SdbUnBUM5C
aebIv7KRM5rS+is3jLYf8pc3lBrB68y/+JdyOy+ngbnAfUuD6PSGT+pk986RSc0LM+z6saoImaaz
Y4Qouv6faQQhBqjA5+NsQbxP1jZS3PgB6BDYNtuNm1mReE4w1qK5hnbMX+bm5w21DsStmTpNHU2+
ukf2FJDtUhoZvG/YFdMM0AW+0037hBPNu6+9YpPtaTgast6FMS9fOX+7ZGmZbHLyWJfmDn/7ejEv
pgIRERZ5hSXwjUR54bmYkQQ8e/3EY7WBH6vxCEWoIEL1f2PYiOg+3aMT0zjKVqDpVJ86oiR4pnjx
pLe57k5XZ5gh3yS4LhgAt8ijhc2zUHPWNyZe88cDUj7aJ54ya7YR4lpIzLJ2PUc3b164zqTt+S6K
aY3+V4FLHgNkyGskB+kjHhjhpUYM89kTfeQRdiZagjhIrcV/fc4IPfpUrC338lSkYPd6uLT1BMRg
x4HHtcV+r/qsZavRJvnKQ8HEPg9A42TkASq4KlFNAx/lh86DSGmmUi9UbQOUebPra+jypZwCbBA0
09RnTGfWjT4QtQL+2eEQ/F6Qig000H/RKxIcgEQieRSJQxtmpz5ApwsGMOfT693FPb7/FT7YB89m
TCImxuS/g9T/IGgbAzHyHx5WNxky9iKr2LfdqcJP0TAYKFva/v/1OFOTAmx7hbsGxvuLBc8s9lU1
GRM/h8SR3A6c6Z0vZ4ehc0h16c9Kxz7rw5N5OinJtjkSOd0oFI1hsU4ICG0Vp0lo51CmsIB9tKID
VBe7EJlDF/+mIZmuYl/ydQZXXTlO7fqv4gLPFYsv1qwTnad2xNpV7gzjLXl0E5Wv6d0IS1KxJVxm
hmqmf/8mjATFw3aKIKDQbHfFbWpAm2qMlcusOKpo5VuvtsCgRb7gEC5tLpI74YXgzzJPN7o1Opxm
DBvdTQqGK4eqyCDh1giHtCEANQCsSYxJo6ttZnmoCXgreIGddXONqoBAe2f/9Awcvk1qWPjdccFD
Hv3XtpWhynCFRVgbYA5EdxNUA5UsFfoLzAQaHxR1evT9GF+Eyp7rPWeu66bzblSmRmExinXMg9jQ
2j3dY5109byTBp3PEl1oeHoXl7RQUNN4an/Sx43az/U+Ld6Es2Dsh+mposAZhO9RRfyf2CjpsUFo
ouJ57Rf0H3w2HYsCh4Gp+oLMXuRdwdhQdndSXtZ0jDk4b/nyuNR+aLI7JvfFLNGbaqqNRgvTi9Km
kVcHv4R0/HRHBK6NSgQg6bOlxfZMKyO2PDi6Yz5OQKX1MH8rS8ou8gss8IcLn3tOCl90aJSTHXYx
XQ+GP2+ZS+14WiR0mopVwplIpg2rt0UK2DguKBBCHN8e3W1vnTq+MjlkHle1qesg2AytFgOKrr0D
AYyXQeE9yeO/WiZzJ6CZtL9OqW/6XtPI3iMwNgEUpImkaRhZMqQMYm++vaqIbKK4vf9lQ/pkZfwR
hHpdn0YzUzcL8sdKgJLsZ7qGl61pXoGwcMf5D0V5NA5uxaBNpnJIZJGE54GCbZj/Qq9/h4OXLAZ3
jpytterDsRBYn99VJYH/aH4Pq6Qa9c/HmCS59GwKeChyg3yL4ZAEKjoYzWmxxGDxDxkm4DTIO13P
7YHTsDtNVimDsGmCykQIU7MR3hJdvoMKnpWPkEWJ7NkErRfJIYUiuw3kzQc+bTErOyiK9bYEVbxO
6rXF/lzQQS5Mt6T0kB9emSd7HArSSzmq2EXd9nrb4xoqke9rLjWe40EkXRVn/XRRKcnEswVPyxiL
+OdqK9O3tgDWaqLvX/kj2cE45S3fG2zZS5/hcLeE56YDjHzCvhWxRWwbpPNycfEWAyHXlokjFZqy
QKlW0S0W78tKANrjeZnpqu/6oFHuQiFO4MDleGBRvdZNtZxb9fYVWMtYDGsP7dE2BSJHvdx6K2PC
75gsLFpiA/LA/RtDhbvHY20+yKGjFhnGpqREv7q/aasmC/c9XEjKEFuNJ1VqtsRAXL672i1ntEC4
2vFz3YJkw37/qyJA14mCPTkTa4nG2jv44oWtX8R0dsXqrxn5/boj3PKASTpeOgAYM2hncF2sFXPf
WEAqZO+XbmhA5Eh7n5Ez3fSIUfc0+fGnRAu9ynJdqf03uo2mKjDeZmGUAVic779yrDP5mOjwkIxG
Fk4peEcy8C1yIic0nRCwlQTWn4wBhTcMnyORutRU0sRQ3+sozXJXzAl4pmQZK1GZfhmVU8kKe6il
hE4VcyatF/blH0oMXTlLeFxF8aveuMhWXwjYotykw3xvHuGX+pzGCtR3HmDBD+puZfqWuo+zJBkh
A6S4+aNgz0zRNzeBWUBAEfAD2zB2kyzweofLYCMdv/j5tNtJIpgBAtL+ft7i08eI8r1uQjLk84gK
Q+ItYBiYRzj1CEF+MeOGFK/A1KQLMqUZP3lUWiVD995HJ8fWFyOx6IFec0zB+WcSpXY8N8IqTG3F
BDYTSXopvQo0+X+cbOwEZ7Tewn0PKmfSf8dV4XQZ2hPfng7BxSG6R5yEnaJl60KonowuHiFwZf1N
GBL4NLWKN0PtGq0mj8pPCYlkGSX2iHctUMtvFwIy5Gn1aDNp3EH6I3hkMqckie+kDdc55xkNgmhY
BnVpXEoClU9YJFrayaL9RMMbJl3YiGF4FzwyQHnGpOYZbXE7zoq/iL29gWwH9zD5S2kAxe2R5rmI
WEL8akL8N3HTBToESRi1TxifFq4yq36fru/zL2Urx24STZi4Z/6vm+xMcC270odbKBlc/Qy4lB6N
GxTIsxbIlKp1FdbTJvLQy1q9DPJ36Ceb9bgZt/2d3i3lDBAL8sDfPMCvKkyNvW+aPsRlOE19MIzr
OLZh1UdRhJhZ3pFsKpjL3CSaTpI89YqKm5bikHdHz33HITm1aItDxgfVyDW13UhqEmhdUO8oCVdy
sATmOBmQK0WkVJ53ydNApTKG/PFkGFxo9welUxonJdPa65xFYqTOHttKByltPKWLUYrDZaJsGGFP
LmkyXRur07AtThKiZp/7pXtA4qgn+20l/GnRskQoW5wtSgP2UWViyBTeAEC9aLvL55Ddv8eR7oHF
OgBOO1/Qsir6ZbXgu3ENkjfGqyY6CO8DaN8pRr3Ch6s04jKOn8DJn/99M3M42p3MD1oRbSbTn5Mx
NqpzrSN7W+tNJB0Sp8VheP92btX6HbntyD87GACbvKaW9HEdU4hudS+aoIsQ/ylBoyv6FCipSVe1
YzalwstGhnt51gUQX9ytL1aC+Txjy+PqQJq4/vm60TD1dQh6tMmuWrMUieN411I17kK/q64o3Ptq
J0luOm6U4XykbU+Sjb0ns5wWB015/J63IocUJACljytDuKXt6W7O+TT45spO2WjsYFTJ7u+v5qn9
sB12HSwePcoq0FbYl2wDoub0MpqTsb+IqLrh3zqxzeoHm5kyuwGrI6p5eidJG8szMi0g7EjobRlc
2YAjJASCuH/fsuanti9QrJH9OjPZfxoRONUvTG+SfTHXoVwhgkJVO21I9zSyrELvN5RbPXHFdRC9
viue8z3kWb7WTKxSjRHXxnvPasyv5pm4q21TeaGXtZpwV2D6NSNorDcqL/o8viE9drq2gn0Xd9y4
uSRrGUOJr4q2Dp3L3WtnJo7BG/oDa34G1TT4x81m0eFhr6nwZkJKlZIyklm8v9Z6XRnim13o9zx5
PLa3PZz+8v7BDKZyj/Ka3JmfpRY5V5oLuEtkZGwKRWInedHAxzZwz61PuGkBcdSZsYHMOqV4IOQl
CfryWopFDvzxr7yTK/aE4DulnozR0Zk+mnpync7m6OomWXYoxDgR/9MdBVHqVZCa6MK+bcKrr7sk
rN7eUZlyqR6eVa4ivN/aJKprnMdhTFraj1KcrtllkCl/c6+OZHaHEmajEkqXt85kek3Chr6/BN20
uJ5t+vmOn3jNqcp0djDTK7ydAZINCHtgw3UZyc8ZybXUALbEZb7TnGiT5wYVKQn152cMtQ9nVvFD
BX3p+iQdtsPcILzHRpe5EI0nBihzEeoCKx4l8mv1Cu6PbBxswGPDRBn6HK9IiZFKAmJtFq/tmNR0
aBhyYIDOdQts58oYyWWmQ9k0mg1f0FXBr/eXLQiSFEIRYZ5AMnw1uzsB8lNkfX30K5oV1Rwd3BYf
r9uRQXG4oFfACYk8iFDqNhUZc7GuJJs5VNU0zy7mY7eQs0bdVw4vPrxS2hsPuYyNF7PY2I/3p9qy
jjA0OyjstqW9cf1ZF22mc9V+9DbsRY/ebrceuxMlaTqkn2nfjsiEqLaajj/cVu2uRUDkZqjlvQrN
oSwxX28wcYK4WVcRXQUkDQP9GyksXhZGfOJZ352hwqBaiqPplxtMf5GTklEL3R/bpeQgQTD6uA2J
C3R/tkquaIGiiVJBQrPodkRe1lnPSSfBjIUo6FqJPNxZ3ALJvbEyJUhCd4HwSmOY5ePZhHo/PK6i
nE2H7F9rckSx03FYDhkYKNvniJKQSWztfv4oEZvp15Onf/QePORD/Iikf5ORLiXH4GtOZ+mBq/GO
VxvMQHt2cglonVGww4ftQ1hPUEmBCkQmws/XkCknhNM3ZsK0h4dWcuu14wW1zQKHT7Mk3QBzBlVc
zAkif2kRUx6YOtABb44hdMGcWhy5+IdCAo48kRet0A9M8LMA+n2xz5fcoB9DKg1UKzzlhypZ3Gbx
8GirNKeiclyrQe3GGOoQgx2r+yvE7pzjcMFqf+y6GR2TYf+sUZygUsohK3mVj5wvsifKuzZTuJD/
sNJjL9TjT8VbaV6Tor8NNcW3HV3IlUsfR2jkk0Fh2S/DbLHGvHEgk4d+qqBqT5uhP3BdaxQyuxFA
HxUxc4qbtieqOUaDKCME+NOGJCmPUMoaifgdOcd1/yhmhkL9jUFnCZB0C+TKjgscMuS6pWe2Vj1d
2bYkzp7VMH1drkNpOQvNGUfmr0skK0MZo/nyJ8n143W3Bpx6dzmkvujyJoSbx73qidV1kIsNo9vv
IZa9V5BtXTJBPnDEXB/wPmOYnVtCsWpewUgvBE8X6i1YrUSSqdvmxbZoOA0/5PZza5IljasVvK1/
4cdxB/fbxKYQd9vCQJ/5Ii2D1OmxDBBM+90rFAhJ2Z1Va2rkrYRUoH+fw+rUPtFCiU+RCVkcXoBo
gd0QcHshum4dfNe79oczHVZU6wrkllNfW3GAGCju4itQl+R2xzN0vNc9G/bIxeaMYuzb5MQc2b8B
1N8/0xmbn6vhDA+/N42Buv2TeEe2OIvsLwfEKaKzY/Jd6EzEq1XJXfXLmvlrWYp1FsH5+u16yjLa
A715+W9axUrWx49NfiAXb3DHtgPY7xcL5kSxfreSL7Kqg0mf1ZCVHzW9GmqFWz+nXMoUbcFmq99J
hJt+42/fnBvIWTjC+MKUrAV3tcZdtRHzxitdKfbGC7rNIjCePX1C7bFpRY9tF54h+QIsmE8GSvbk
tQyiuT+W7p8mgrro0PE0pXIMwValDGmkEAtyqUHgQgdQbE/VgIDcTx9T0fMUp6rsXxB0vT+uLQzr
WL6RDmAw1EUTzM1J4UIdozWOmZ+ZyEjAJWJcF4G3Y/VYkTK0ZI5WZhFzPwKYtvuZ8gEzR9cgDDFz
MwbxdEQMmlMJBeQ8aJpeI7aN87ap7o0HJx/SKCRO7+ZE0z5BW781S21GRlNUZFo7LNzW4avD1Zij
4j4SPvfgSeIsWBQR6pWTkQXkP++wUGIHZQRVhEyyhKc5VlmdCD0WjPFnnSY1HWAYh4xPEVnaU2Ev
jeXpR+jz6RajbXn3qcMWJaHnLZnL+DOhZ6QPtFxVjvtINA8Canm7kGAOaokrk8JgxmEJxEaVBjk3
34iGcC/L6kuraGSdHc9vS7J2XF/dU2u8N7p7obs0HqOu7zO+H0d05JHxPlRzOSbI8815phvjneCW
qEphF0GS6qdDCa13FftPDVllGWXv/lfjrF36xReoutDRNJXa1kwT1ewjpULQu3VMJsFitKcfQezR
LgQAF3GFpgwPa9/GVKRnsaTJV3UmRSUvuE8oJsniE4/SxFoWCLMBVL5h2m4ZMKLEnmfGE77sO6Nu
LTaeTVhSYiZqpqArjJ+3UwFTTzeXOJUFBubwJnd1FeO83OYHeXMEshZ0surcwhHgnLr2s7vUYWNJ
1M56Zamb8q9SHFRdE0AB01IAbn5CXKbCgX23HaRHvIseljPDTgqG0z4ohW8qnrCd2hkFdf3eJJ69
0TmXhsaSHjniKqd3TnDEdhG2LT/Kh3M3ZHci9PHGcRHV4UGmeHW4QV8zV8he2as1sH5EP6PI8P+X
Y/K/v+hlGivxC8xXmuGT8m9PdZ8K7TrXnHXA6zGTWs2jlK1uCrCREpJBcRaMBWg6bA8fn793CwVD
r7vVyfrnFqvTVnopyoAZ1Hbipd25s6O1j77hul+N7/c+sFyDT6sHVptb95EOS92Yz9saRZXwbKI7
nF+P3N631AOlrZeHUJmuwm3XrVIAbHq6ZjJyg1YviyFxVqD0IVcluUxJD/IGp8EYNrRxD07/QqrT
e9bxLBQ+aSD5E5YAbq0khCnuQdTPG+ZTR9FR5KJC9Rktw+J3OiRKdFXkC9bcIQ5AvlI7xXlwjNrU
BR2z1IPfqYkKzOOoxREdx256ZkpNtSyrUU4m8MaZupuXiIhX9HIYYpys7qrh1Uh8f+v13F9TwSHx
gsY887lQKQehpCRc7qzwcX4Bdjgab4we76QOUWzrY39Dxr25uvdAr7rEZ3iU8wncdR2JBVsWTl5m
C45guQggvq0WBuF5cid0nYWlU8+85dwPBErNYDRHSDsrXg0enTXj2ERZj7BnAGwHNBwEdUZ/hP94
X5CeZppI2ke4FI4hQ5tAhUZ8QUM2hI7hzRbMZ7SFAFtH4e+4HixGRCuNC6tjwD7ZOKCB9C5Jal+Y
4WxZyJjY8ZW+ZZwTYlPZipGsePksAhVASfeoD3mb8I0Ntf8U2ha4woR/gKF7zkRzOklSCv4MADTP
j2+A8MF8FwgjraiJWC7GyJ6wWyKg8ke6qXEMHK5Hx7ATzONH+JeOELttWVlztNU0oYVpDSXTIMXP
EEmLEmlDXcUytWBH6E3TVOTULweiDnt5csY92oz6BP8YJITwg6YZg2AYrwSnDvx1mGNY+b+mzDFb
eOQOjlouUxMYsVFPl2UIi/4Vdt2PB788m+OWrjaGcwusPE5UJaalc545s/94K/PwFDGRbMG1JrJU
bRtjkSmpr+AAyo0+koM6lCjLJoRtrOGFxcns+zBrehgCzgnpeMDrLqnPAJ5EB5xLdaJ4zXzijUnt
CPS82JbOtiSei8+LO40UA1ivE+wN0jQIrhb5f9Hyxt+mIJOhXcA5mE/Wf5rUIRZNCSChzypZGaWG
soOp2g9oav6Vq/qkF2Xyt9tuovtTpyi+2Wb5YHLnJa2VUb89suDqmgVk3W1KWwoxcGBkrbLPb2YF
20xckQUw8Q5mZzsgzRfacmNZnq7kopCcc9BRUKSawBnM+QKnqL4gDY0OClYSS0cMoylH/1aomNFO
QhTfKPxXeXSCnCyg6xzFn2OcZ/sxDzxZCkjgfNPjBdbiOltzeGi4vD6qeX2HbEFs8pvDlYx9kCPp
cnKo7cJ+QB4n/GaGDq72FEI2Z2UZzL2i6iJ2NunqFT09g8/RzT2grV48Lm2ZzeRprPr6fEGZdw8x
Xc86YatflqX2p5ZzNyP0aFbPeZ8yDxH02sXcOixKNQiRTKIFWULS2nfhTCUnrCEAUc24M0evZZXp
xk1wgVtMrQWZs3jh9iS7bFlL8os8PZOkPaijEqDDYo5+e3Ps0+DxNZ3AcxAesPrGE9f12JiPoDAm
cPe6/4Fc8jnRTibxbqQXEppaACCOWcStRpMl+ONcrYMGYeYRBPvWOB2lyjqia0HkA1Fj0UMqMSLv
CoFSsYRNt3UoP9eE3kxuM8DLPiWcPsgHK9vyvmoMSyxJyLLlk8jGQgLg4sO3/njA3wiN+JxFo5ju
f9KHqMZpH0m7GvJiiOqWPgpzJ/f4on3vBxJ/Jjx10Y1xDIT8jnpoYeELJZRq3gvkn3wkugJi5j73
PyPbgiItQpco8EphJPnmferFO91gsdbdl2LrXguQhxLXQUMVOpOa/0Z6wyXlZXkp5S1MHlvEL8dR
E16htLaxLGNVRbxhLAUFJ2sIYSgHFc8jMyIHzZv+NHKP2r/nTP9IdDLMaoapxF8vl9RtPLFh4dms
KF0tPk22D2Wi5KqqA9gUzwk4KgjO0a3M+ocK/EG1UaiokKEGpIK0A/GWlUVrY++7iOlRRv4Wq5u+
KKvik7wipSDrAKSqM36H4XbK6EpfIunj63Vj6XshlX+kpsbxpJlLMaI+2JbQ6BsDLIyebrcenSWY
fn17hVFuuQlRh9LyVTbK/e0P40MXPEowl5uqOyPGNd2JRUpWhJ737XHbQu01S5WggzHPBOid9pCO
QqXLw1RPUrDLSHcvlX6+sM08nNjR7QTs8zYtHXuFyUe8+Npa57FjlKE4D7GhiGEoqV5vKcNjU8pw
9UurcYabacB7szGIQ2CQN2ngHgQ6hgN52Nytihegk1/5Hq/qi06xRtxEpwDsIiEsoPBt2H57x4Yo
VNlm0dhhugMu1sNU02nJcPcso8KnWvmPuXbsHGwN7bQMz8PhPBGBxUVGD76wXftXSlrs5s/RYi7H
6zH75O++Y2H6eVcURL1H3IIE7dj5ALtrV7t1yFgs36hQWycSK3BUY4ZKnJewCF2EqUqnAH0l8hIU
uDLTONuS61flKDZjhqbhmjtF8LJhqSuwLrobS5KM+BAW87A7thtY52uEetC/v/+0bb+xeqjfy2WP
oWv3A/6FuuoUnjkP6ZNdzYWcToSHHEinS0YiDn0BrFGZRH2EJc/U9IH/khfgT06Irb55E9Cw1ryI
UVaVMzts1W6Qo8IvAezqHvbH6plpTOx/CcPIQyRQ4FaE5XgKb2J+ifFsDjH6AJnZ55mfLGIELLB4
mH6LB23O43nVK3wWAMkR5cop+bwhjpcJ+1q0HOxZ402o+LM9VGmRSoKcicEAzknsWP0XpIc8I1jI
fHuvV3wlE/M1tDpCmdxClUDz9Sd6xlwFPWZtbD6BfwVMj55LYpvo9BtemI2PzXqGXVDZ9p+zIXdE
GsbknWvA8DgMqixG+hsKNjqjG1vYQ4wrZgiPH0+FkAypK76KR9jmCCRj0vMju4FFH7dTuPoqGP3I
PS68WhNO3ojSaZM1oUYODiTfHJoWUAfm1Gmf+Wy/0se7RMbqhUgtSMyxC5satnu2sP3EEvl5dFdL
/tAqRn9G+4HFR4+vzv9uzdbu4/V9+/h2Vj4Qgcqq2ghCCXRvw2nxJvkTF98zvMnnZsiARPJ1uno2
RamF2goiLeDDXW9JI3F57pl9tIm4RLHsAzTa3oTuOpNIMYl4QFZiVvtRbyTKXUoWICyfUzo+4wTJ
6zaDPnDGi88JHcPRAlKhmsh21/FIb1KtL3sGXv5nA9LCMM18XiT9zWyL4psBkseDcpNHrEimONqI
7Zt8AiB6kP3cdk2d8I2zXCLNyVZWvq3DARyq4109cDStX4nrUWn9eUVQ8uHzbqu8ufou9obwXHNQ
pzzJlZ8iKK/v6z2C27lLFoKh3rTFjWrDhujGaTFQDOO3D4V4EaxD6VAFoBbG1fso150kcIjop1WV
LZ0WmUgwYzQF3cWCvYUy1JNxUEZ4Pt+9gEuElHwch8+a3hDuMPr1g59Mpi+xTc9FCkA5niad2CfC
v53UOd6MdBO2iTxKLALtl31CPJpVWBDrka6NLUv7aou/0DEfiuTBcJ3QbrbzjGqZTgDZJPKh4TDq
qnbPtsATDEpU3W4ZX/kvWV2eGUkvOP4nULnlIPLsART52ByS7yIQqStXes9s/QGtfO+MtjOLtFmW
0D5hvCJGvi16QZrLKFLdlFPn00/yxGN3Me16BZx0d6kjr3TOITf0CkeMA22o1mTqV0VaulUe0PHD
8vbeUm6hAAfBZgOMzDT0pZVhAUMlkeywsIr2Pc0kxAib6+Ooe7DbKoPkJGd8qYBW8jiL4MZZKJAh
XQ+9qpLhpKMr3dt3EWjlsHOxVoDiyTbuz23Kvs88q75VJzrCW5xfPn4S5VCxgOoh+nmv5gd3U5IN
EL4DoNA/Rx4MlhcFQbUQ+RRd0VWKxtystOFYd00m7hylwp1WcCGqZtHDLc9hKCfL4WZUrLqDEdAi
iGiRq77TgoxBEmbCbXfB7WAXg966xKosONHglzOHEKBRxmmIqKfjVAsKskTIJG0ey9lmxYmrVaGo
RLc9IdpmRiBlwg7QWEV0S3vn2Evr0ywIpkhYc7+D8wk/X4jsg+kqJCionTpN3CrRivJ1oGM17Mmy
DZiq+5VtMbnlBnKtN93nWb3Heg4C7kxoFBFnh6qf0NkOZCQyHPq26apnsExrVRdbzFN5PqoFPB50
R7LPGDvUHvRxGkrghVBEsYquwv9O9N8J+2RQ8DMO6uiQfUMsTK0Bcb5MQS+ppuyHpIOxS/LQ1WWs
ykdhx4gWnWJ2HC6lInasWI37i6iyrN9zF3toLyvMrgKVQfKOGhBsiXI0qULEBbtsa4hgRrvhBaFM
fomG9lOSXUVtIe3MpxIo7acsF71CFwZ/qjau3o52Dk7n76/3qlMSfZbG/iLGF/UyDcMeQzpERp40
MCIRNt/SQ42h/UoGSoG0yC0pv9Ui+DWvJ29vfhzLea+YGfdToJStOov1rcGpmOnxWUm5hWTPeUTy
XO98TsJRO7ibWjUIiyLSBxvI6gWPsZ3AJK+VETyLs1d6OzMUZvnY0qgpWm2o9zdU6BduRbLKnE9B
UdfZLRNjTOv5J4KlCxoREL1sVuE2EVy3JD/q7rXhBwN00yjO59Ea/Cez2ml/m6Z/ilGBluCgEFpK
meLQxiDZcBWM8+9wVCDvRSgHU6OwBdwfZRNAX2QcOg7Ed+nzSn+5qYkXLtnBsjb2lDhVcDGXwSK2
M+BcuJjJLw87fREHq8yAvLGBrtY/+Dfm1wLXAWSNzJ2TzQ16QAd3BaPxeObwXrXNFUTWSCTJojie
b+Pa6/+Ws0RFjpVpxarcnkHxmhBvnvjnURBZztP8hkEvHtfnG1gsvfO60u2wl1YJqE5dlNffhqnJ
Np5zrpCqW9dMkPCxn9ZGuN+LNiIfAEBSlpn8MaZRg08fyE5XVfs3wcI1cDFra48yru7+cm5xTMPP
3HsHqmsxAks4yuEj0jObxfZQfAdg8y6zv6bOGWwm/U3K8ae8l6avRcuI3fCPY5olffg9E8ULcy4l
vh51PJt0lbfHOAYEeyChPIwSXj8P0PfcMED/vJWvC+gfxurdSJAnoTaDELglSNbTc+DNy/3vEzxZ
YxJDi8nAL+fuS0zAYaf6bdvZDCN+uEaR+qyAc6FYI8NvQHFYiwj9cDzIlKX7ki0nKgAa3j8QrAdB
UDas/rfDY5XsFW0a+IBHU6SLb8OJIcs06cjEzaCp1u515eAidE01NIYLV+ArOhJ/KnK2QKJnzaOK
wbgDKWqt9kp+ojYqhhjaMAHAt14T0hk2mGr+6YuMS5A+c6cFGd/x+/RQI6L02LvNvGsX/NhBMA2n
OGB7S1utuC+K5RlNY+PDKfQkACqQyruCf8F3/wQUCYW7ff1vnVBXCM7bXAoDH+xBBpaOs0hDJ2u9
Xvgjw3KONzsj2kZ9F39esekSv1RL5rbc+osZ36N6COEX+LbAj6W1Ueu4OqFgI/9/7vielKMCgy9w
tZ/+p2iK/Hid2VGuZGUybYkmsCFWYkv7b9h+hgGydGwy8Kjs9AXJChdzSESbay9Hwag1pyr/wMPd
V71aSFG3nfHF3OT4GQ29ooRHhSxylzx3HmGnCqUFWjOupZoK6rQAkPCsYhBnwk1WDAGD8i36J9Pa
ctUZrzM5EErq0WFhcdkAe3kh/hbpcf1Jf64aMahGCVt4SoNwgJXa7K7nVFA/Wks7uiF0BepW+iy3
nw8iFdpEH/znLW8zKArGGwvUU9R+Jr8pyN9Bx0k4TtnLRj6GS0KGxlrKU7n2ixl7WLmYi37XHooE
YAG+sDYFwa3kqnwDcaCLFjG3SxsilFqe2O0VmjZGKC4uv3ny01DQv+CmC4Atj1x05/y2ugbNGXhe
fmoS+vAHx95C2bzCn7hcPomPu7APUDkE8ZNwsKORJ0PQtNhAATVz3mfYFoH9wQ96NDiqHKfwRL+e
VXjfEbrSQGlcZ1WLyztTCTvrF7Yrn5UGhx6lGlqZDpTK5yUCcTCVfa7+dG/iC1pdTrEyyv9cZnSa
tmlDLXM8D2FOnGmiuvgjuh63SIgvW6IrGMwTOd7etWhPjC8PkMNqAjAEZOYqYEeH6Af4XPWPBnVc
jVFFmV5FVt6o8TQyNzx8L+McxleyX0uM9I2637PRLGXRRvVJ1UHXluMYFjRsb7ES5qsSKtvcDKIm
LrwroVt6psH7s2MPPKCltpP4Z/gBTk3gO4v72TET+af4T02nywvjQh/5/S3cWVqjgoeSVCM7vtFf
w7YSfXFabu0iD/m+baRAg2Is1lt+r8IOnJTdjCMuTICs4QnaRN4a1mZWe8G/MhCnBsgbCBbbBImt
L5l6LxMNpPMxxZfuBkyyqTLIL55LnJT9roXI5mvJdeagKWi089Cz0EZ+9VSN+0n1/MF3SfcjLEsF
xUcIYK7EmwPza6ydOlMt/FgkAISSWZRi8ERjUMWm9ymK7pLUtaEnoiKYPsebjjYA9cqhupQ+hI4L
dT1zJpL2g+hJqB2pzSkjQiDbIQm3O+q/9GE1Y+R03mzsedt12y5l5/uxHXcXR9qSGNIHgJSKGzRV
rOhkWduwxwilvEp+LuN5w323nv95dJgR//V97C83kKU7zsyN98stmCg03SkYrOH959EGC8stbsLi
lLaqFmLGyANjiRXw9Z282+73wbxjQYg6+N7Xz/WQyFXzKzmyNRfB7+HnlK434ip1iyXrxDVB9BLy
AO0+tmyPB/XCWjeE7IVGkD3DMpmVtcrypjdPcV22YDvPCDrox10o+UN86gKR84Tug/3y0NBH7Uv1
h8nmtjsXuCoWYhTG1prfTPLKMK/qF0RF+DWXSuttNcScRyAbP8tkb4HQcwxKTAvcQKN8Qnf/E2um
DZpCdzLtDQ3IW+87mr+6jMRVOJbiEa/iYtPLujMeoxRXwSvRVhW82F/p12uA/5574y68v0Tb+xvM
s5TsEuRkFENYds53XhNu+uTiyZRRTe/lWGc0ei9xVGiRHbYbz0IxAPAmZc15ZZUd7dOtA2m5TI1R
hI90rPcIqNd2EdrHvsV5oKaiDxNK4FfJnY5sXOvWYyFTpxClJTt/kX5tThkQnm2T3aql1BSFHPXc
u/dNsa2FxmqD2jVViokpWz9KeAWJxNRcJlrtV5Zu63Pa4mhalQH0hgodRg0y+zVS3nDccDCOTMJ2
Jt9JFmyD9dhNQjnVESq1OpjLqKqkql19bVwhjyhB4zNls5QvhB3LoaGOI/F1dYU4RmsbfIuw3rPp
QMx1TORUFJHsNvwIuKGG4jPOSY4CeQCucqW+FF/f3q47WCLKitst0ZfVBY6m6ppjKRK/oaEUWZAS
EKXZyMa1XlvS6/gRuXPc0uRL/26Dov6N+bo7CoSiWqZcxFI5Ol26drV4mze1pSijNQPLt2uNCPwI
nXLgnSctkhsF+aqe+rZfvZRT8fCzT29lAMVQwqJSFrMy4xL0y6nm4eW49BgxxsCAPBLGPVkNHya1
x3sGsFuLqZ725DHTM99Msj236C5QCXQlZ87BP48JUsZ7jkVY32dvvTntKtpNdHKMEFqUtKMXBOCJ
C4x6/s+6e8luv3hSvUpPqEs4TJ+4xOsNnDEm3uH3WS8E3b+7aSb62I68dz2mMEhg9pEto63qinyr
kiCDJrXj2nxjG18IIGSyUrVsG5rLeS80BJwwrEEFTZhVjV3Bfq+ZtvldGtmJG3ndMafl0yVpKCQN
tv1tfzt9HpEFz5Ma6TFpIwy3uEA7BypwXyCtBKcuFBp+8cyHHdd3NnQ6nFT0EHWgrCSh0vU0Gd7r
EK6S460wfcSCFU2c/YWdNZN01LCZ5jgQL4bWYvWCY+ymOg/gvLoUFdCZ/pR01fRnYKcrzO/udKX4
40bUPrIsYoarsW2UqJ1qM+VZawbUsylhtI/BLxvkPwQybsd092NB95v99ESQfsbpFYUmZZ0DaQW2
Mou1kATpSVkUF/CqMiAFmQvctjdnn3oGOqcnnNO0AdE+2mQfWyeT86lSe5a6Iff3y5e/jHhOUpBG
ND4SYHOgGxKXUl0ZX0aPbSs/qgb1uCs8eXb3ALELowlbT0KOM/xqAVuUmFavcF+kuwT5+nlDiBij
TU298sRrguWyC3hhpPNkGxixrSXIj9Kp+aWOwSqDn0147HagxVY8thqm4yG4K9IOpo9jnVIk+Uqp
2Bcj1as6OwInqLrlfdD/VnDSKcjhGBoxBtQEMbu4+jRKJv1EpSJoGBEhXnBPc16GpZcPC4h67sWE
3jCRjsuraI4jLfU2DGn2Zt1mmRo4lJQZpRoTlwTUBl3cGD5rZul9+z+2/wMQoPkGPKVm1GD4T9mQ
sSA2AhVaK4bnlybmlTpJV7UW400gNgCCIAlhVLFuNU+qWBKH1JTIl+dYeS1O5tNQlIY4D8IbfDIb
FYzeMphE+1elWarXmXXiKviJdmkF/rEC5iTJ8XdkDHSzH7lgoEMagdjWMaAqmSH1cQx3L6FDF2LT
BMF4yDOB2oNQg0+vocutIzzyHjuJSxTxFNvcQtfjJD8ygNKHNGSdBaNx/SplhKxpMpLW+6+aKaBR
658TF9ZbaPh2MO331X6aiHmJNoaE41xCNmjPODxMNX5JmqI/+28Wlf58rNJbwARvITT4diMvrfrd
/xVF2Lz8XMVN7IlktfOHTeeUwqWUn4qbcE/Y9OR3PjGjdVFdYLZSbqhhxURPLf85EdKAiX/aAoiF
YF6uuf+7D/QZLjy4Cnjr00OObZMtIk1bp+yfcWMA/ctIUU+ciYfzPlzafCpTzbB+TYCMWZIobGei
wTMN4I1OeGuku23aedRXqcd4NwIclMjDzDnaBRTL15yQmFM1KGFiuI99Z/6W99fR0stoMQZAhd76
Mxvwze9IABFIr+gUbi3lqJPw/rQFpoU49Sq5XVoOrRfORCHpYOgol4xvcxrv9tSaKvMIhWNtv+dT
3ESchUkX+TRx/F4CsWC6alYSOY/kMEQvlf7rLfhkEOP1yGZQM2hWxPEYhehR5uvdReqOoJiWvhpD
j/fLAHrPyqFA6q/JRPezupNWPzPv+0XtU4WTPNCdBXE9VPaFgdFtLTHJv/SzK6MZti+72j5CIwww
kimRdMf93kmg99wwryr5FNAhi20QePmogyuoOi9X6EGaQ+wsFErKdmLhSMJ822cA8wz1FRfCGDJq
oaHINqU9ygIeaV7FDoGwagI9VGkvhOoONAbssQTAITA2n2FU47z8mVdSs+14qYo6EqMJlM4W93WS
H2aDbM3l/n9Gb/A7Oep/23rmsloLDWFmD3SSMHcNqcbZl3Oau6hmbV9hwww/RqOFaS/ijK5RKscQ
ojQxB/0TQhTlh38dwl2kjBstBW16a7QwiFnPlW2nqXM+FQJR8nLZ92aOdQMqkvwU/QJN3SwZ2EUw
p+nOUX32koQPdqTZULNcuqV1tj6GTT6DnxZM8K1iOf5i8/iIgk1Ndg0MRTplF2ApPDhhFCATGKkU
h/h9D/htgyIS8YTtz26Pdl2jl/8ZFmTu98Oiiurp5AlgPg5IyNSp5vUbbpEe27TkKO76ygy75xZB
5WpSgRoWqRUTi6Sg9kCQe95QID345QinS3K5lRWu7XA9iOMFNsPpIyEIAylnffRQ55+3JuvyuKdy
INHvGCnWhPjb16yilYyUCFtG7LTezMd9le8cqy/ZCC/FyvnpaLoYtkPKnfAVXu/kBFvq6fjeYxVP
T0bgKU7tUbOuGK06yZ4EwzJ8l4tYX9fAgUfcRM0eiMFzh/YVRidwD3QH4486C86qHyVqzCBnzCcj
6/WH0euTxHbXUXQBbsLavml73UjHtMj4EukCF7Z7u27/wpZZlbvZx70ai5fq2yULUHxihoo7aTac
l39n4yKEp5xbBmAVx6KFoiEXmCTuxlIvIEGxPEQQJ1G8LqjawLuH2Dbc9BN77n/CiXVAWfyavb7Q
mx9jEsiUfQGyV/6C5DablWQ0DB/qdu6XJF6OuyKAHzHTURrq97lZu3mVikCwoH5I01hwhQcXTIRe
dnGVLORIlD1UwlxL/ug31+L43+0XL98xoeQTbluCX9rLdeg0jU7F4fOmONIV2f0vc+eNN8N2AP/k
WlZ9G/7+abvP1qwLYdoJX4UPqzg3GcHMB0xuSmq1fTmjNHxOfel4UVfsGsS1OkWNsxyc+dzcKYXG
VU4J2SfTQWbbbs+SlnfZXUKMsgBR1flDjuLE+3dij7G/EZsWaB2IxpdkWdzkIDFvyJ+qCHUIuLKE
JEkF6Y7UFrjzJoeUSQUKm3DrqSwdnFKkQUaISc1ImTjzpe1Ezz7lCn54uW/VfO1dk8kFzWwC6rDN
GS+HA+y6tAd7UBA3IlvzpIsAmelPmPFZSC8Z8vJbaGzLSLgZpS5ezLBfK2PIfgK/AFOdO+KCrdks
xtELkCj+6s9t8bd7ZGtulXvRL7Z3fDvI34Rb8T8bAYO8re3dLCB+USdbf40DNpO3yXaAlnwss6xH
5EmxvAJbfBK/U3e/kyTSKT0Uvy0I2c+nGVgk8jN3q1bgZqRkBtcbW1P9oikpWi8DCP6WTiHgF+pY
xk9SO3Ip6CynoZx3Ivrg2EUWznCXQZPcv/nCS95F3prSBN0QzuYaViIMbEDk74syflGSN1WnlAeD
RqpHZBPocnN1qb8AnA2GN7i/32S3NfL9g8DfdXR2OgFlm/Ye9bvdvUF7U/38/lrQW20h+b2nxl/d
HZPmPjwKJm54RMDDygH6AeKfbqL7w/3WYTV58hQEOu6+imgqO1TK0QLdsG1ykvC5Nsi03Eq/md8q
n1Mp2FQ/IM9/hy74hURccjwXRUTEdghY2hpQWSpYBZXIR0eKk6fTtHI/yLIZRSnW9tvbodTTVp+r
exB/oRGaLyNCscjh4obm1G77OyBi7mczUfS4M03t7icM86S5esDahjD4xOWHr1JLCV6lVqn4og6e
UEbaukDbBCTiMQPIRuTVtafTsYreP0uAaD8wWIdWw4E4EV96VG0dRHEOisY+2QWkpilmtGst1P9r
L985tNRcQfpkuzfjy9wZ8uxirjsAUsU1dlSfYwizfZCYqlVaKKNyjd6OQLsXlL3dG1BMvDfIGGLj
ZHLZgIjvWz/g4V9RlVn68M9auCgV2LE7ERBj/0jRM354Uk7qNk8xPHcRvqwWUhBWGI52J1ZVwlGA
ONAxWcO4n//D8QJtff1OBpp8H7BxO3mxQYelYB1l79MbWbgdCTl2XdQWHDDvpOCcCTk/RWc8VjHF
wWE83rJ9DMoN3vvlgWyhHsc5UZFdHpUYIIjD8a4Y99Khls11jiO7qMpCmAQ2uLDCHnKqUd/0qT/F
cszWbg8+o1pubD4WAA3fc8c+2wsDtndtJUXQ7UrL7sJKF87AgVtBXSxEXo+JrPqlSogplC+WM/c9
ikmU6wMsbckhcvJupwjlzGBDadZMoWSCQedLf4X6SQKaMtRNGkB/Zb8OTcnCzW5wfcxuGlmqPVC/
UHBWDvzp2Nfj9roLAWj0rPKZQkhVTMa2BAola5fkHLjNFa9PwfqTxlYY5rUz5lMixE81FBQQal/n
Gtz7i7kfi8BAzhTZq02giO4a8RPif5Xfe86nyhXKJsj05zwxVMtrNCEwcOO0o38YeStU82gzeAPo
C9MJYfQyz377Pk//E9wYX0gNwebTcMdXx5PJSINhps2lLLvEz9U8d3KfvksjY8ruPgx0S8MKLek3
VmmHoiV/SWFSrLwQLcSfqkimhpijiNTZhpOXZsziMRSqoQgx7VHbQ3drjYgHhrgu7D6n3vRu/YeB
jsfrw1QYNgX8nKvGwA6zxEOkxpExzXnFiOmz0Q0rwTROtERx6ZVFOS4b/m3tGWWoJCgADAWnNbjD
pED8InT4nFTyxwB5mmDwE6fky93J5C9iBjUPpGDh3UI8eUz2KW/OgtHjaILqLufyn77w0gaYtlXS
jlyc18tZVtUE4kbvkExrgMA0Lbiz3bIemIXwxixwKzgxpxC4X4aZlHlFe45M9BamJd1AxVwftGng
axwuwoQ0XWSUDrhIkCYy/r+DakJahp5sQiPmyH4xBKoVf9dnCFAIBGP0hlugy7ykCpcQC2wzM8bf
bVZQ15u3vqP9NJJeUFyON07vbR2bKrphwVRbAQeFNbGvz65XbAS/IbFU1IQBVI+6LWwPic+wzylo
WJr8EGLekPI5NhI2xRMEsdCNE3myAPi1wqezoDmasjdP0c7L9az6iUse/+5D3nBq6nrc4iuw6rPQ
k4B1MdVKaIkFpn5sZNHX1IbpQgVCl07o48ItUV0YQAkWM6JDADAL3z38wvT3UsfStOqTTE5shYqz
QWdEUH6u84uLtU5KXprTwIjEaDvYfKWQvaL4Cfr14BxuJXhM92Ni9USnZTl5WvAbHA8q/qy2y76p
DltWNoKOmnxbuRGAaxeP4HZWVCcxzCPr1LUttGw4ZGBOCfxoq2i20LzjDMkQ8oNH1i2Xli4fwhJn
0kaFurRCLymUPIZZdmbSlTa/EWSVfxIOHmSXXplMmAMiMimNHJgprkOnykEv4R0ue9KPAQTatd9B
wYHLGte9kwq6HZ8hdPhGfVrpSTAoU246lwZ3fwMn/NmeC7X2SlPQcFdqYIzLjIIah+IBimVWOTki
AtACFbWpIdd2Bnpc5YsH/Rju7Jx1ouz6yrrUJQ1evcqr/fSlEV06kXX+j9DDL+Sa76UIRaCyvDrW
9Qnx/NSgOxW3sXVWb4/fkwTfjoohxG4vhamBw9x0XRFrVOi9yGTkxzBtaBxnc27lrsZqe+d5jMi6
44AAIJ2T1AwTsqNcbUlpY4/8KwfEFUO2JdHyJ0ysebUFPqLqxROJ/dQps/DfkhaZc2oFVRG75hEw
X0phpmsehD9q7jXFimVssQPLDO1GoNU1wdyIOCuUVpyjNFI1ZOgEfN+0jjI3T9XPSokujELB4dfo
HYFKjfL/sW6ZvVXJ7QkD7jOtCNDlsqUCWDBNLCtjR9ys4dKG2XQcCowjQD4fz/GqnPy+9ESD/wZX
of0Bx6jHUgSShz5DBQMs2qn3Lk6C/l3kOjE3Mb+Ytb82PQPKsxyE+/LZWzkvuAeO5Hct0y3nfWI+
m39Y8TKw8SzsyZwInv23x8UDYzWGlEMC4BA4mKaRr6japRkCre7JLnsvIWFUyoAnpV3XmbTpupIX
aosbUz9w6oqKpq3aj+Iq65YdtynnqYIQTLH1Ac5DVOKuXx/bJCR3FF8PSBlvh8Hl51ZxQjjV9FnV
L6ZoUmGzuqPIgRa/JGObxcM8pCiJb5i9Sfp9J+RsRzm++5vbwXeUVadWtpBe6zpR0B0rBo0lf+7b
Y+6Xwlqwq1xpPRcAxY6I7pwU3NwwXsQM+fizerSW5mH254htYN0LyfPBESbBgWEE/iXOi0D6G1PL
jrghjhSFDKx3F0LS7bToYiWE+M9CicrLjeMIONaVtg0TzC4j3SYJG93iu3NE233g3dkHxgepcAgr
bzecPj3HDcrd0eN2OfUXhVCgmhZMPDQL3ppV2daqMO+seftIczI3/6fKVwCSAWuyorO4WMBSt9eI
8bpv+GoHPcrmXAq3rT2dCrMdu0KEAZweTWzjeMHjJnXZxr2xSRUTClDe6QRh/p1HXtgtombZWDRW
DN/NCPqcNLJw9NV9qzArF/LRqX5xtXkLMW77a1iOIehwQU3D0hnSRtGNRIDQUnUYine+6Z7iJbBu
wC5N5SUGzP5ObSdYD25ykaOtpjN2D1Jqj+9UrjDkhH0dMBN2EAcSg2TOV5k3QJ7fBRUrgZLUVe6+
cClA+VrsauoQfME+eJbIgBWtC/4V0X3ptkLN6R76RsGEs0YHLhx3434gxwcw3XJgHzmCXfUiUgdl
5FjdpZU8giB4nammv//Qk1RkehqNWrkIZpFPQ9vnFEQiPOmkz7PiyCrKfDYSATf9L++53aDjrCPW
xuffT6LM0p3OrtQxr89FRqbbR3mfPBnENAgl80cF6jbiEiM1LDoEcSflR99Z9ZJEr4ARQAZmb3JO
NzXTI6+a8qMv9q87pMRUdqd5zmeiBRNYKSWcJ8KN1nd9xrwdYyBDYFV1IctFDGPIf7B1abu7W3xZ
6G3940pBJJDOHF+2HozRYGRQv0MLpFTLtXZgrv3ixEh771aHseMBZk77sF+eLT63c/SyaLsLRzN7
4/vNioTt/J+yiffxjgMN6OJRW/vcDqr/5m9TWDZo2CAIALdo7QJHj1DmYGle+rlsg8boFkG88Knt
ZHx5BlJtzCfSRSeLnE4JBhgpdjXOpaK/cGMzARhMfnbKvE3vz7RoYutUdrpdeOJ2OOXO1v0VVcVa
ZA+3jKxDHi8N1bxxDw3pOYJS7J/3FZBSR0kOOjvg1zZYQs4j8wRQBivxh3dKDi8K7t16Ni2hnt25
Ce6ZtZsvgRYzEfPO7v4K5cQD3Ti8xTqlZNRPAOrXowoi3cynVdcd6fwtfXI+SwLF+PmI1DlnZfj7
yARO49gIf2Exe1j6cwiBA57JBup8DQBat3bHxjru2JiZKcrjlEfhDKUh67WOfx+sUibRApiow1kt
YESuZ14jF8S5u8Kj6jW0OIAI8hfmsKyX/kt0DHfSfUBWYFvR1F6a06X4hQygbPWcM3PQehTMNAiI
d6Zism2YxXdiIZD8p6Jm+ngfi+V7opIMZpb+GMiwpFHJ3MjiM24fiKzacZdL5LMgHLay9pyKc4vQ
EB+Xsnql923OAazRFkS+7Z4i6OcSho3GMgPU2btCVEuRMrdWmEiL2lT9Mdb2OIVQ93DeKLnkRJDR
HPRtMqdxbw4n+ckDDFcf+fB2tQn9sLh6p1Eq672GTn+A+hWPyK0PGAGDI99cOFGDwrrKOk1i096O
DnPOzFmvoYkv4yoleBeyEgnd2n3GsjWbWSCAqc7LdoDUEj9H2vrYY3zZ+od3NwJuw15M8qEeVIOL
Eo99K7Fq91DvJX47CUrioWklCWv1nj6JyhOQWBrhB6XNXruu7KTHMIeT9MN8ai5KrFwHBNkBFJI9
Xh8rtq+JsZRBznnbBoGts0utG0fMtf5RmtM2b8sF1XHuDwEqRNgwTSQSe0HHAzUbRSsrw77tdHst
aoG/XJ8vhfm1blEaHBV7WafC4L16N7i7I/zYAbHpyH8UmEFtDDnPGz1/+izFVVaC7wxZuX+Z2/fI
G/b/SmNXa1IOXHXuDPPRc8Yk/F7WT5AvCw+J7ZD4gEwpDXRLFyOocgDdOv7ip4xQeNTCxL0lV6tM
Ra0G7w1jMAflklTC8I2nFXUBt2lzkESYvVx8A+5BWALM0KScR8yDmHsxsM9SWvNasCD/19Tk/wy0
hPRO6K9U8G8Kzlm2erDT9SR6UNODi0abMrNiStktFRYyRZm4Mu8XHxmikiuYfixZg3XXJ0IEeLAJ
Q99eePNtwCAuPOWs79aq7dyqjUV8W59YbnISe8+aQeHAFvJlDvuLUgQT6xKyf5iyI5xr/NFuwg8L
ENcKaN1D6q617oAIxY4wgWhWQ4Y56DBQrK2txQnLCSARqZ72xzaEfCEUKjpshYwLq7G4kDSmvgJZ
2ZLQ+zUHVp5YS97o840872sV1elki0mHNZ00EnhpL7KpUqcwyKAWPTRhC1IUgiEjG0HM+Wa2bZbH
3+Zegxf4N3QTS51cYo/WqKJEFxmZL3rIUsc+EW5T+XYqlLW+inxOThCyhBuV586SBekE5q8LGRUT
G/CzbysxkBR3NxKxCObLKmB7bJwZvv08El7/6sFu2FT0N51/CFQuwlJ2ZVeGW9E+1VwGq1zVRVyC
TpDJ5JhPEirbpsUYgnWs7c9vWADyQ0VSdY6qTRXlCtEVmtV+OnRK2WTOaIb7Ax2irR5hrqK+5nXy
/sVoZUtoxto6xj+Ji2cHCelREkyHNWi+7GOohYk+dkDKyyoVvBLyvP0DheHqH+4l6MIJDUQF65D+
CadZyWQ06b4mWG/xD6NO5lLfBnoOE8cxSrxerJMoR1okhFG35CKDlZY+K79nqvIKrzJ9klR4t9el
SPCdqS0QCZN+ZpnR4VlTm4uxk6bHypHx2HNdkZdSVnGi0BPktBowNzfGD9u7Av/4V5btJ02MbyaD
ULJW1QNT8k5a3Kf0OcLzCpgO06+kZXvMkE/fnP0hZ/+rCs8YAvU7/jhZbzBnSuQS3Cho0FS/uIS6
wOZ2LRooL3o4D3FAtSblym0v5iFaR7dSf37ZEnYl0okcMtT2Mnu7qXW9sKlFES/EM/I3wsoVdtAl
2N9Q1UjBkjooMHr/Cjt8WCCdiAEU4Ov6QgGNAWWq2d/mtBcjmAweH03dd41e9K5IpvvXBydYtKDA
qjpwezJQ6iZan867FCf3Jy1djoRfTnZXJ/EaUIl7UtW8N5BG0V3leeL5FzzBw55Q+Hp+zW+eHvBY
B8XneFNeLhjSP06YlpACBJR7hX6osjxvQvUOjMRUXihg/n9RGePp9S2RpGROI60LUfg20+etP0Z/
41sscegqUzK/5PCMhN+yRzlG71KmhwuquwNeVdUjnIQq3fhij4LMLY1sf1OoGVD4sUICOkY0EVS1
JljMfjaNwPk6/flgdaDjfi6r9jZp/BNkBU/wE8Mis93zmiAjiHG8w1yOjY8XWhIWXcwaXGbUe+aQ
kN3l2jGVCacRtz65DlAv5Z34ZNKMBhezBAevpJS0SNNZRUw4EOtoa3Ch/XtumjhmSCuv/JHCKcqG
hoq+T7SWFejmq2RCLjOc3WoGH+1fOd9YEtU4qu70i/tTPVkOWEzqBxv82Vrw/N84hoPBb8Ap5hZJ
YZtgba1lEwwmf5rYZ/YeATsduqYtqWRMHYrsaqFqme1OPQX15OpvsZxNMQG5PKv91rF57FoyV7xC
/cikTueQFUezJJ7MEMYOYBv5Lf+I4KODTi8gaQwMMVbTOfN0UfnzMc+myvrrVx31NLRzH8kkVTi+
50H5GwOFk1nvdS7x7Tc237bMqt4oc0QwV8iyGTCMLL5xWkZI0BLE4i25EFpFAbuAThRswJQels1j
oIGnDHo0AG8/XH2lmMVGzQ0P5evrKgsdCA21V51pTuS2hF+O3gWH0xKZQbLzHF1EGlTKt8HQJmM0
ifMB6c9oxRBZUJ+lE9Z1KRElt4zYZp4GiiTnAlT2+vDa8crJbphVeDvCdT5+TBJf3erjzGmMSQiu
WFYEWm/xa3vBq5RVSD5yw5MSCaxuWIWf0Nm9PFiu3FYxhCVkagZ1N2vxZjAc0nt2XfEg3buLinPR
jtQjnYJjDz4ybVk6CeDB8zZl0F7+wSEDu6d+5p+T2Pxjy0NuL/YuMddHmwbZAduQ53EnfZni7MwN
BeISvss1aAlU/JlZ0pzf/33OEjJQ1dqcc2K0bCjZPLuEkWCq3tifvxysBAK5VPRiMmVKXJTFmkUD
0ewQA3GbJg1s7Z1JGAXm0MdQnlkA0vQvnvJZ1LfiqQY3UccpoyMscDmC302St5xLlRSViefZUefJ
STjiK0nbW7qlSvtNDnUQPdn/BRch4Tmp/PPpEMy7ms/xzVuIAFEsJC13EL9denkpNqVXSocyxJuI
TUeY8vgWeXi1qWMQFdPKHK9LDIWjhz/XXT85WbvvJVqMJV4cxDa30N4mYfL+HqUcdXv6Ka6RloLt
bNijms3wqbGnMEhk0GlKzsRJwvHVksQ1OaaarXWA03L6bwZoEhQg53uk2UFIvEB26EHc1AKHLYzr
NiIpP0uyvzL9MmbgDN/iMplRpE/lTKspkKSNvm+wgopuqolStIV7bGDHhlpm7eNOqRXRPfVNZ9Y6
KoBEPNIoHDecuNwV9u/8rTY5aHIG1/I/EIt/Fm4X1biXgKdGpa8PjRKO7/E2aLjavBfTmTrzuEfN
ZAC2jfIAhpi8UhaM5O6zx7jmmfRQs2KENVrritrmi0QlloAGp2FhE9hfky0EqN7XjIGwEiQxjVrZ
RNZm/q+Htf7iahBH3KLb1hidrTv87EQ1PGJWG48vZ+iNDRj3CP6tIU0lFl9rzrHe3e2A/Nr95mI6
AvrcpINP42fIUSoWZmq7DnLy4y9JtbwNQP8O3yiObNZw47k/YrK+hZS79IOAAY/CVAqzDe/P4U8G
PVz1zPi4uFgl4CPjKX0uWWBE5WBZhGGCiM/dbR5+JnUKaB9YUSP/rQ+4/FCnOGCNiJdiQXsEAk4t
veyxJMr95MvBRq0tCWvYeW7B3rqHRXyhVhHgRpkMBK7iHi2XiCvR6MD1oXcR2JVB/K3DCa9NhbKU
Isja/zWlw4MB7UtB1GLbAeZV5A0RQwv+uS2Yomt91vjjjz2tyfKb4aVJ7qJtE3PJa4Fx0gs9pfOj
hM83N6cVbiSqPBw4xJtkhdpF2jBF6QMOBzr+bjOGznoxROBkUEYbDF4j9RXKYTceRk+rNAbzdtqM
2eqpz56+4X/MPcEpJhiFe94AY2bR2iBFnRoKkxaR3hwclahqooo6ypc7/gIKt0om4lvb1dLCqmDa
gwf790o/DuUXE/XZfLc6r+4E6jQNqyqMexyC6jag0z9KVChSGNQ2j+d90ZxnP5+GarMNc8AGczi/
bhW456tO96CSRTbVhLh5g6cR9ILQN0rld/s83mFbovP98s5whNnZIuw52AyoRtZEouhOJXezl0A1
5yaFA05WEuuV2Bxj1yg0Wql5WiLPfX1UuGdx5abt7qctF+seZK3fEL6aeRbMA2dcOCGeJd5KUlrO
cS8lLVjkHxRSdACl0vuRknubAXa2CdUojoYFf5QH5WeDviIpLlMxoPBW9dVTywG2weyv+JeiCcZ/
IpHR/74+I/A0z0jSqyjwrdZkzM0kDXj1CJWEZQ14AZCVEzoS68xRI1yq9SAaZiIfVvwKqlcfHgGy
iTtciC+OLdNDtSF0NFPtGxcigtP/+Xcn011VrmRpjXKvsXer04OmWBtvp6BfTN3hrGo9WhsvWFPI
+RU8JHJi62ProX6n9dIxDpFzLaq9X6cBRsyYAFg1mI99Q/Lfb68iHO6/X8evsmDRDTGeWNB6Z0tI
OxXEalE/2bc/47A1kTxuIn0uASrRm50cbnJS9GMKKAWPbER3vskjUdDFkL1z2hjjL1wjKmZ+FEIL
APmkDDdi4YCtynaLF7YvGepSZcH2NXshQMjQr6C70kNAh0m4z/7PP5EFexJoYSW2N04ODtrbhl9G
TTtB7DN9uG+HwF3OChqfYnLrYU1OsCptxtMDryNKSUpKvC2ZQGyldxOG+DHUfVeKxLyOIaGtQXxM
ONrwCmy2JNJn6SUtRxNFCKPS9M9zEYo/NtQJQKZiJ3u5hRx/4zc1J9Z3d7/81yNuqEzZ944+63Jc
iYOGPVcJndTv8nlqfrwn9/KtodiPBQBLVIWN5M1+1hAuNO0RQe+mE3OIQdnx0oBPey7xM3mAUKxE
S6Vsam1kCmXWorhyjxBPs7nfxbxF+rAvmenT63AXHAMpMTu0TqjqycEnkG0BSidlgmP7lyLNke5S
TeNaPHGjOf0Sx7B0rrMp4oZ1Iwnwgtcef1SGsNQ2W6tvUseQjbhc+ud6qndZkGBNYKA67/LFKln5
P1tqgnoO2rn6lFOi235RmEoL8egwXqryY94BUX16ZS8lwbqIQkp+UUSt0SvJAkrCVb+8rEQWCJc7
xZww479RVpB2H9Z5bY8fQNeXmlLw8r2Oc358v3DtrXBoeCrgtpcFIGDkXgji6oyXBtOnTxK8i6fi
ETVXRuHfKk8LQGavF7h0gMebOHitPpUjxfzxhoYdNkP57WpAX27pGXMgN/uJlQSMxNlKQlBhUIkQ
qkAUCSmd3J4hLW9tNY/PMF6buzD9VEk4Rd7KqI2xslVvh5A7IIXCOa4L+/bPCCpOtxAXk5irfFYZ
r59eKvF6kbI01sDcTk66eIRFeycQq5A38g1IhsU/F9B2kwpgV2ZePatQv93o69HHeg3K5WeaA/WB
P/vWWJcyiYA5373ASVt7kbPCyaYya3ZLFL47i+zY5My01CfSr29Y/lPWn21qpF4GC1NvdOh+3d59
x80VNcte8JxsdK7pd7ZtouYpXfIxAMRHUXu+F4teyG330xctH0QQmM/xlMjCzmo9uaB43yMlHN0X
CZqIyh1aMGVEAdhinWz23NxmFxmgZlhqPCkhKIIJnf5TKCEQnzALxNYf4MAaUVh/ytpfO9NHRIOj
h6qYV+K+zxy66C2++3TmS+ZwvcRDjvOQUWDzm2RqMWCA+mJgOUT9VJvUP/Mq8WQWRtYM/SD920UL
SO0tS3b2DGX6Qhki15RTGbEnCabZmu51LhtETA+nWNBbI0WaXf7AY8wQAMb7Bs1F2NBEB8FgQ3an
Z1eIYK372g7Vwkoqpza0yUdFKn9h22p/1y0cJB0RYkSd5fQqEX6eSxRgIlH9Ylxc0v/gRQOHSnhg
yLSimgEX7U6kOAE8qteIP0cJSs1PavoHlA2kbt92NH7M3myHshlT1plVLlqw2285SEGky8PACwDl
Vf6jTSa4YSFXWGMkNOyANWiwVhnK0Gl3LHp3M8iLTwDOAG9L8+2we2NBl9rIGKbPWIVkwxQX4DS4
Vve0Llx41GwaXrNic5lgtiypzOc36IwGUUbl1ppRHzD0qDfPuwTgqEbps/7pEQOaJfUpo+kYRAOh
k0Vs0MykAHoNQPVri0AdlFZ9nurTnlcuuzFrc7m27MbSOQtA/bRvXyc9OUEI2b44Q59TClX2GQ56
tzG+JL0yKuN+mDvyQaJ9ElVKU3b9a8ANRNsR4bTEbZqMq2tpd4nw0G19VjHIBukEPJinjUIfJNii
iAO1G6LkZHMT1hc02ahF4XK4hQCYe05g/3IPURn/WcVcH5s2ZhUpROluY4MrrpNy+TkglDceA2Iz
bu8v2mDsig5PQrhvWQm73tghpY2qC2OPUylf6UtB1WAr2LiAUjSa3oey7sE/N9OKyDkZBew0ITru
5nnaq1T/nG5LLk2kkinsn0jDabLbEyOpqqIaue8YbJquXEFCTK5sWkvpo5Xl4yfkgRe3zuKVPiqd
PsJm+GD/JuULp0f21/nIhOmB/cvz4RaNJx56DoTy6r1wJeDPkyqDLz7n/zBwOQdHQoayjAHFZsZm
T1O8iuNK79dhCGveRkeTuTUTJHTGctdVxLbRFgKtOBV7YySCPDYUsqCxggBInaEi7dg9audRF3nw
HZ3X+EZuJAbstjckWeHvtIYuVSJQ/kMv9fnoUvBmTQGCm7UgvDYoPUVuSL2gmNM5AwocZv8pfGmU
6bE1qlVDgNboYf7Jyj3QAwzI3/4DOq7S5M+Dzj8cnQcw+53fiCgGdvfldCDOWHtqiNnYQuR/9kXa
Z8z7pPJukDuEsCKqH2jaK4fxUbdq43Z5ZilETEoaK2d9YG5yimIOFzNgvzCacawArrnYUSN+jSRG
fDwwlyxVCBTbGyItv2vFFxZltZZGYPoOo+jm1Van4raW2fTwn9KE90fgj3pDouiVaDmiDuVrBwNd
WdWFAH4rrKB+d1M0IX2A8rucGXGQxGNnxMP+se1eEdrde8WTHBIq4h2DZhG4EVABbaqVQIqE44xM
4OsRxKb63mSBbRrWZxa+rxax5D4eH1lOJ0oHdYKlTMQL+4oSgX4ufzGFtromEuoszHicZAYYeDv1
FjJtBYcpgLO3Smk80I/YG8O0R7oHjh63EZ+9JHyxGzrRKBIJJjujDd9Q6FlZD3ErtQHtb0J519R9
K1rat6MJCNZhEoIT19w+KBB5vFE7jdWlEVO17+aZjuXsikIW/u6WnQQ+tzBeGo56ycSm0Um1DnSg
J7c6xmRSSU3te5YsDrHksn1Kh1KI09rNCwpSPE0pZtRrYFevYdmS2xhn/beHggv4zpbG3fCsyqa8
w3nCSkCzrLcMcDsrkBYVGuHl0sdK8A9twxbBgRYHuKx8q/mc7OJ/EHwWfbpVvKxj3VAkRX8aJRs0
ePP7gOhBkEcf9TKoZlJDIqFTDIAsVHUlb9BaAWFiamplL7RmRFqJCvV2aqzF7MIpJkrPnCt/mIV7
vUEwg/1eW+5h1dLuWGpOgZL1TW+uQ4gUIv2a5OAeuCJdUa9sgRpodA21pk4uF6NksNPC1SmvlUeP
gS+4UO0x/lJIvO9P7grMrvF6CzOZ6p+4SQpfQZJSSCWwjDyFozYRi4EZiVYCXahSDzFI1DjJBahp
u6UFCeY3JtJB2Q6zIb7rrYPXaC/HPa9/Jj81PEagKE9T8ASt+D/en3GgTjPovDtbkmBy7XBDpDu8
Jwi2p36F9TrR34b+260SnzIldnLBlhQ8JaEWNmYYNs+N1lQLaWsEgwDBIn9yLyZkbaxne77eD3MF
GFpeuDNnxn330htvVJtp8k24VARkEBauq1/AeztvP7ugFoK25vcP62T4ay5CsmXQuFwCHc43Aey8
3OL61slGjPtIXG2PswTet8ZlpK8kLsZ6kPfxs3a3Dr6e3Cb+XVe+jJ7f5gAtOo5owmYxmf8RU2QV
ZHKXM7ZqIWnnlrlXsE0i+/Xyg3mVjGzqKGhjHf61LOl9IU68JzyunjSdP08XPMGBB+lNwBR+SK77
4tklE2G95AM5CRHjgOU3ipVARAAIu8UftvJ4I29if24rDQCC8sAqYasc8fihnTNPYGK0FpxTvSdU
qHzbGvuKds+AZ2uUXO/FQY3877hsfJrpzO9WfrtZZe5XAD+tvh2oPdTInsvpbWxYvY7PbGqMIibc
FqYR8/XgH+xM/w9piB+SSIRpb2T825RhlcsfHHtlDWOjVc3OPBufqgxxZy2kWLtjQw55EbAXPZQT
xdwHbWhRgoFq5EvBjhwzPx3kLm7wgQdsDZhWqw8+5deCIljqnlSnvIMGbi4MAI2DS8v3CUEQmg1Q
Pzcm/DxlREi2ky0ST/M/LK+y3b0hgkxw5C8o1jlQvu0nNBP4a7xBur2H5fEPzQtwin2yoYSbt+Kg
Yt12u1kO6J3auFQlmd06VlZ6o7tNNCobaer44Wq809Dzr/BCYSCB6bN46zrPYaQ1FDXULbGjp6Mb
qSzUwGebuc+damaJ/5g8deDV/vZiXRfohKfdHNhlspZF5UJd5vNU7GEMFUa0ddmTWxeLTCtNQzEU
3KN6DVlfRrTqc4Pr9te18ea2dvlNYC2mfrVtnUosm7lhQQs9cuPWs2hUDJ3DiQlJMfXQ+rwKPKVf
PUBAhfh+93UTuKGz1t1vHAdwGlA2ubcattypRDr3VgHAxqMf6MHa0mQwkWdktJMhG42FXhLhAhB2
hAE1u/nCrqc4iJXjycAYdA3XqZ9VMmAy2KvnPeP1VRN/UGmsLVK7Nmk6eEHEptpIWpAGEtu9qcQs
hNa6mD4wFFluaDy73ezzllY/9wOyzoBDxTDM52aIqKxfQauOt8R5fBZNOM0HsEpHchESJxDXUXin
uRplBf5BsGAnF4ynJ/4u142VE8XHtG85vMHCWccVaCgYJ9jfeVWzh39GJSRxSgnPKGcR5ETCP3C6
/Dnns3talZwQh0ZpZ4dgGSJvTWlfTuhnO6z8FWZBOqAjNBSLjB3RM9E7EPk99yI6AZ02wrXiMI8+
Tmp6tguzrpYXQwPA/QLWxvzHTKc6AzWOwC7tC3ytaE5Nq1KH9FrmvYIXd/q/W9gTZFzb3KLZIvtK
KVCOBToUt1pw/kuK+4qdD/VzgWdLc7xHP53Tke8b2eg+sQux+79kxAGWOXuQLxOs637CCXdwuoFQ
02pdmfQBsCfeuwr/L8HMG0Oluj9+P4BVARvUb4jiU2Nq3/+Tu6V92s6U1FlMP5hN3+z1luu/kHaB
xIqLIT5U/tMtCN4IodK3S01v9liLiwDFP8qKWuQo0mx+3tiwMOM8FPsXfq0L953fykE1IYUbVFxd
exmemfh5pOaK/OG4LkuSQi3KeLbIOSKIEAZVFCocfJHmuelcy3pz+iq8+ScP8p5T5jBlOAEA5PYK
5+HwiR4Ut2rB5MXuCyEaUOTwX9GzusX/AfBzvFYrQY5nUmGidmH+huD3TAQ11UC204doas87hHLA
xeNxrwGTkRS9Qw/HHaFi4urSdSL05q9Juk/ZNk0fkfnKaXnqjKm7UugMtpNJkgIgpFiWm/pROpdZ
nYEF/lifNd3Rb+GYAe4OyAa8cqw73fS4781F931/PkLHaXlYln1DEVDCrpV5PkCwMQsFu9hOHlDV
DiultKPBTRqmMMeGbMpc3+eBT7RhpFmxYSvhzB8ON3KWnPxPncCRLzELDAzIMleA9tovkdocMEFA
U2fTGqiPDDgXrvAr8/zacHOjyiOqOgSoeHQ1Vo9uirtsSaFKbUu+2g4BaHsK+zJ6VPw1ZIQKbOJm
Q1QQsu6fw0lw+5JA1oxkqF+L1ppHy/Lf8eIMpVEVuhPgQo8gFE4JHYuUnFGWgbd2MJcuzTbWKCqO
7jIscainj05BWhDSn0F42ZQcNB2eRSCyQOsjPQsp869XJ8GVCkCf26zOdHt/opBnWd5T/NkAFbub
87MLvnmv7gg8eh9X4dAwU0KKpkizFS2ZFKrhoWoCX29xl5L2IYVdZLo0DRRfnZO0GN59rao0BV56
NXik1FClicvEN3zMbMgPhlIH6gfJAAbdcjcBm9cooIRDXMVCJl5BE7jxQcEXGwKY39Hs8Lpa67Y7
ScUH+x2YbXQCjoYbqN+nDHl2qRrkelxYXZjWuOej1n/vRlCPMfhETR6eb2tivZopC/1Y6mJTH0KW
U9vb6cTtNxkVgVMC6TNpFvIZS3FehoQvKPFBRg1mx3vmHHOvfBGh/4HaWsXMKHlmIPMjSTApqYoD
Q8ipcyq4CyV6F7o9PCEN2hfZ1887V2Ls3AUKOgitoXtSo73Y90lep8R1nlmJ773Qt5NsG9yWJknQ
zqxM9T4w9yPb4Fyx82wIe15j3KB9llO2WovqvtkFJ8rk5owS+KL1EFvywVhk2h+lwlzqogmU1NS9
0yV6wIgEdW4WK03TnQUGs9xDlaa2JySH9GglNjtNgOPvWjeFsbiThRoUrZikxy3hlv7Xi9cGqQNY
vWZRSwiSccOrK2g0foaAIodgJ6QLBKpuuC3uxfwYS3ggdCsx9P5c54JLx1nLklr7jxKETcLmvjo7
N4q+L/ULPFidhaVTPOrj4Go4e+E/R73ZOznK36N8AvXNKm8ku/T8jOdgKk3kI872Q18SIxYp9qiP
eA1iyxiV2K7gVrjxIJem5QwQ7FQB2+wnYY1Jhg68NDqKvPj3ciiuH4YjQ4KDDOFmcGOvEfNFWlxs
dToMZKwqIAhnw5Ac6c65wJ7qluGLK+j2p0DOj7DM9J72GhV/xJbGZdO4MUB5tuh2THdOvOHKO0dK
W/MNXbvpAuxb1SEBwQ7+j1WfRaj7xYElC4aLel/PVgUI3uYWun/U77JN6mFp88ktYUb2o97QtPKE
UHayiSDNgQTYoDg9PYv0JZwL1e7TY0FU9GSWcdio7CdMLSKK6GlOVeFMMXQHK1mFGoqw1e9/+4KD
c6eMzgLK97xY/+EUl6EE+NvdrF/PaYQah5U09+vCwgMhVsdvkWDRVzFGSuKwe5rDpPR0RLEolwd/
xueMKYB+nNmf6v3hWWgPo6wF+tNWl69CkR5c+/gAD4qx9ClxAazYtAHCGzmjFWCK3UuPW53Sz8Qr
BVvZykKNRXdz9R9ldLdDorkMgcZ0XvtDQxUrg5rFiPbU6xDQXtOEQQMvOqDn9B/YgpOGc10zC6mo
6WF0Xr00fDM8g2QXK2fD7g5iBsupZPvC6GL6U7mwcZBAUdO6MP+2szglCL4edOqXzVTO2Xre9bON
EJrSgaizGQtObYXnRpu/zQKYSvg9os3+zZNvHWO0z4aXpfWG2ypHxbkdA0ZkgwwS/j2nPc32Btvh
SaXjjuDBra6/QVUetQvU7kGnmRdRS9Zw5Bn5En/TMPt0outWIUO4ONEZh4kCpNRdR+C5Mad9/Jiv
FulV69j2NubLH18GBtw2hP73yviVKYvdSvwdx5TAS3AH0ZJC6df1W+tR3xd6emf5UjZO/XrGoVMi
CCQa61HqZ61h7ukHEo9ietNLdEZXbch1qWTrrMvWxqMTuPTiCeyO7FcxSS3VBFR1egKoc+qaJyUl
h/aj5tas7Tn9ETrKJV6ODckgkBgfJDLI07EmeQGUaZs/Y31I3fiwDZgk3JE51WzEXAF4WGCGuNY6
1lJPjvBaqYQ0oaET8em/1fnArfiiMe0etUC/ja5LH9HV5gy+WDoORQMa9cwPp7X/kEJEZk4XmT5M
lWniS8tS9vN3AANvZtWG7j3D+jjTWsMuHxxgi1ydJijDWJVFB/V8PV4Qvi3Glkj4Iy4mTXWqX6UG
C1robIYIR/7gM1JKkxUg2F/L4y+puOHHRwevOBaOy8qcNc3oOieLqpbgXfbIkrA1+bCvD1iKgqQF
DpXZ/cBcAeu3yGFj/WmrN7MV2egXB81cD4fJVz/Z0CATwZvo1YYKTOht23BkNWpNCqmq1VWTqGvZ
sbAlVuHpXtoZnElYNMNICD40AYHWxp8dMmRTNdaIpSe2be/zyiNRN2fahufdCzrVORLnaYdiJ18d
HcMYCH5coSJaIFQ+D5TrbS2HYidq/q1zh2fFD6F2chffCMEsKeHNtWKS68itgzUI2vKDYW1jb9Ks
AE44miCx6IanHbL4FUNcAa8nwWDM0fabopvNEPeLgiO1oehRZq0LsIWP4GYjJm4/KTbXSzCPMxNr
vLPaFMKBv0m3drM/ozChrXP0sbl0Fsd8U6bzBYJ7N0Hs0IJEudNiV9IMSSiRlS7vaLrB9g3MZ4rZ
9i6gl8cGQ2j9/mRSV3MieZkUpe0aUq6O7xcgX2EpMND9MkZxb9Yvcyv/1dq+z+434gfj9TCaMciw
IahzWem1HYVxECDk18tAxDM+0zsrydEB9gD+qNkyZ26WZkEFU43ZPZv/dimHP8ZVUmbwBlr8BycB
+UXGuPOfeYo6JTKik2MPmO7G/CqQGAatVquB2s8pxn1RyGSuSNvZqqBkrbBPxgXpisf5IcY7Ih7c
ABtNVK5AkjVXo3bcy95WikVvjrIZtT27hvypy6Ell5fyJ3r/0PeQOx3HeEH25YcXNQc84UfC7hn0
Lq7FITE/70sn28U1ApvPn7me6Tsc9P1eu0J2Mc33Ans+kwfesDA3zd+PqrAFK/G+VhzHMIocnDag
bFGyJtLJ0qaW4mJQWbej3FuX5OJleBQsrBVwx9LyIst1ZS2AcYH4TENOA3Ya/XNTQe6DPgvKAsaS
kUl3opmVqDZSLardBf0faqCQ0UGFzMc/OpIqqaoXfM2DhVl9f0wNPiJwnUrAUlelQ6XnAkv41r2f
3JhikVOvZokXLTdsU0VjJ+o8wPG2CN/J8Vs2j9pbjTYFCrJGb5GLIpGJAEODUyTjf8NfRty/c+Hv
Dv2RqAjirIVBk4yUhZS11UaxLVX3UmtGlU7pkyvW4EvrRY2Q7RRed4qaszHnBpytzyDx7IO1igLk
7OEMtAGez2fXJwbl3qxmI4A5u1B9BPU7GrxDdNGjKvC7c4qsWQEhvftDdkc6x1eb1196EpNhZHPD
solf9OJkakEYkPpowGMdD0AKf5nA2G86jn7iWZkPPvbKDeTv+KuaAGdTo8wjczbVxzVghNFVlUMz
KlvB7BMeoIxvgdfDXRcUmXMxw+eQtFlosflBWcxaVFxfcsytoujnLRJWAZMXBXJ9i3HUr6XMi0jd
DysLfogT9IeaPLK+UQduscf2yILrqp/0ves6/q+wvx43bleRvrVTh4O9qkwIEVHZ2GwoGlBbGhVB
0IVPviDicpJN3gB10dHGTnOLZtjSzTFc+Vkq9g4WtdLqMoHVCjC+hCnSpa+kEjTQXXT8R4uQlDpj
p5XgGYGjFeOcrxb3cc244d5UPpI5WM0O5TKPItTItpFG3QiocPvQ8mgHYFbRSxc9TDlDLkVjpO/i
+hX0foz4GREn0ZBHFSDqPB6NJXUetpS1lBPmT5jSu8zsH2VmX1TRE84eLNdafh1cxE4KqQZA77/2
zcw94Ms0mcVu10LTsdIzXZFtQNyjKDJNem1lfYB9LXklb3DgwWeBErymux1lqcfwWK+iA4ATkinH
KdqBfXtb/l3y2/rVjd2mWJP1ASukmzkSDpO96JhPStv3fWAlZaNoLOjZTZIbYU5W8Y5es7Bsvrua
vSk/oktuyBm71SFzRpIM5dqGBLlJFfGVlv0C+Pxpd7YIQEkwRniS+P6CzS/fR3w254HDWApJ5HmX
3U/1jNq6OrgYlGaEbHJDCFkc0bgtytmUodDSen78x0A4zoMPMyCC2W+ZAMnTxDZtbPoliEzqv/cK
YK0AXzaYRnYSub3wgjLIQMc0cFK241bqWO3JYya38GMWz6RAlCp221oIIFg23QBWOoyeeOyxWq1X
L6RkqrJ9+FwUQseMNke8OupytvsQHpTt8Va21tS5yhnYtf+rEWlv8aeaWeKvhJjFBldy5TrJz1SF
SAvhXk0vCOoSwnXE32UoO7DzbG2KcKgtfz5K0hlvHypIyjaDWZYB3EwDzLZu+H2yH9CPswIsUsXX
Anywjwf3excbO18FkNAc5mQXQx1qHhF9mBB2DET6FQeD9SUkHnZKSm1nDUsL2JFl4KzXzrwfrp4E
FA5jzXPOakQHkWNJwjsaeNdkto6S25pnMXHnRYz7Tic6Qe271gIZcw6mred7P5QVmK7iNI9PX/oY
MspKK8ht/Rm0/k367/uWIu17CcFMb0Y+lIb/lIs7UkSXlDp6s/ZnKhKpJR+AVNSDJCUl+EqerJVX
fWT06IR+548taCTsO2zIoRcXCkzQ4AsqANJXQrlGBrCdiScfSRD34lj9C8md60GTVv/O+YRI+p4B
5u5+fSp5Ui10X4QefFQJhe0iIQUZ0G4jHr/X1dfkv57n5ioeEzONleCj4iVKlEJozBLNDAnJdsnF
14ewTA0s1nZ1rtkRyTRYH+gXPvtmdW3vMH2sEYtI/9WGN6cRVSUQakYHSrwRyq5JAhdBC7NePIPI
XRKgkBqJq31u1NHsKm9O1u7Psa0/7cEMbIKbKkuD4NkvSlzsUapAiF0idxF3qui+XAru9ZY7GN99
lwiqfuhGFPA/30c7Wub6maDswYxmRrc+qB/MlW1LnM8g6cKDZDi+Z1c3+4UMjf1pTA0ax9SSj5A/
OyYZiDgv2p0WjAAWynExWwqeT+B4u3EOrL4Ou32ifFssaKdgXKaqAKZVwZZDf9BbF6NLE04BdXRy
XrHwuok2qyUqv7H9j+7JwKNJO5Ti8vvdHiWp3lEJb4A62Mq3N0DFDi2YnUi7DzTfBhS+uXDYLXtc
CF8Dkz1iJv0Jy/tKTKEDElzuVCFSDRz3/XwSQppjJZ5QhQsZV9xTw/E3x/pwh+xhakIlOCgt0vbd
cim2na9OT/MD8mSgayXa/1IqVloZ5rbWNILehbk60O0779n27L5uGC0bEQULMBK/yUrbfY/iuLkm
XFaQW0tPXoFsQENz5TXD2xTdOoe9qbBnaPeQBySuNLVffypsAkUGL5uGmDDrrO2LRX9hVGvRQW7E
BY8uRHDsPs8paKuq3xO8tMYcMpurZNTr3tNKOeCAinfmrHjDJOOuZBsgyhjQM6eCdJ6V4w+mknn9
Fyg0jf3NA8w37g1Bhio/QvD5w9S+/WN+aj88hDTfOxmWwKrx96k53a3XLF4XwYIE/S4+dMQtNygy
IfkoRu6RUdIy1wegFYiphzm6xWwOIc6cIGSnBdOUwabdHSl9iJcDTTh+XWowLTTRHzVhlRr7CkE/
F1I7vI2GEwy0m/TuuGQTz2/nt8SM2j95w2RKg8xFMOsaQHH0qXUBH/FD1av97TPtYWEfDyXe+nqu
7V2yNKjnonDPqaIaaiu6lzG4zN/BRynyx8UYH9yc2pFYijraI5xfS9IyV4Hs2KHcZyFeYrX33NHs
3yt7UuuIzydUvCR6im8KMsZab/SiawbCoJ2CTd+UJvRDw+r+b3oDXafRuy4M2oJmJltlD2Su0RZ+
LSV+DECi8id6PKXN652lRU2Do9NDdVrY8fHoyz0+8Jkc4CuwgeToEMyEdZd97+klthp7YeG1Qnmu
j2bZshkqJ59HtknuVA4MO+mNSj3jXMFkYh6lIku7k1mZ1DZ+II/qRsYekH/6tP92AZCcMThn4Hb8
2UVWO9Iqc1heIWNlJ6fjdEC5EJbu4/gohGpM4XVh9GGUCegKzL7EPP5cpgLUzCkoZ/4SFdtjJmuB
sohiHUIflWDp+Rng9buGEUl5vFynkaxPDetEwkLKc9ut8KtlpL/dMVKFYqkLTXemosSfPGvLvBPw
wakuljNjpZ0fXeIXHLpL10A1zFK3yppr8Z3e8MN3WOhNIalzQ8AhbuPbZd3GdPdpnwJdRax4ZyuE
mQM5inGkIlA1hfZaGWnqC5v4Tj//re68wzPMFyyPV5sDLOswYteXsCjOXW4rcX98OHYSCBbeQ2Dn
u0ypYKxjFsZKaCePjf846Pi2IBg8iFJItrCn628PQ0YLQ6FtyUW5vVKBFucVsm5gHLqsML/vHDFX
60L30mJSnjaRVLBL7gtoBsTiXQZBgP9JFjhgzVE2jLKuW9IMlj1seVdE0i2MqP6Isgtm44He3eU0
yzm8V9fyG+hHSJU2HWn3ERHOP8tmNKN9jUzhXEs3v+oYkfltSQk1OF/sE69o08TP3zF36giacUel
BQHHpPW72o3yIeSwOre8S7NSHfr1Xwk4KaQTCL3CXf4i4psiO0Mmi4ovrkuFV1PqJ1YpdA6WBJK/
hjnrhMRgurg1L8btn/X7qS5oU5zTw8nG/DC4iiqxQWxiSwda8b0v8mAGVYlraQLBWQVJ+ve1l6VL
ZiFk58EKYFe9royDk3qT/l1QWRqsRU0W10mEWuLE0kbQP6ihPcFbKUd3bdnrG3Ai3fRGQGAK+zdx
GMxoASkQ+9zPJVHrsVdCs+Fc4ImtIFJ1OyMCsacnY63PxGZCnZUff+1ZzlPKQSnIICtPDzXSPXu+
u2AK64jjw1PJO+/e/2dzQNAz6n+0QPVCnhq6n8uUEDf7S79/PBhNitPxvde0iU6LRM+gJYDIUAue
5tXS/bVOyDisvUetdHGE3u2VJwcxZM1K6vHd0oPssgMLILFfc4jtqG38/4RSBtinPlBIHDQ3Fw7Y
F8PRu+4/uqgOUYXEj7kgsgjQ08P4pvikFXhuvc5fQ1XnkU5gnrQ9IFxBvjp0EK/AcC57cClG+HGE
rr9QUyeyRpyvi22qFRAmAGzkDGcF0sT44JAfv4V1h5QVRwq/RhIFEtLz2XD5icxFb983zvBPEJlF
FPBDuN08dntbeF0fywRg0pNDQwzRCXM43XIWVj2GjJEZpuyRLKtFIDYu7q9cHFabyaZuatfzI+1z
ezeHKjJ8KYNzmszY5uHWZDdGPQSumRnymItq+vyRFWWs/5FGxVYEamuC3IwsYcetgyu3ftfizoxN
0tCx6buQsq0a2sDh3NYHIclPDoNlSBaUeu/UfBemgPYJ+S1NBbxvnm17rOLs11S4dmrbPDI70kqf
8m5WgQW7e6MNKkDIjF86uCzQTva8TBjTeAfKei6/WFbH9iKeUf7DA6X0RpDL6/j8ulImEgsJf4Rl
hnKw/p2lTxipkjIODMyz/Kzhd5K9t6zUWUAGSwCoyHgvszIS+FYwhMvModh60Q98QDwPWwuyBUTG
upyvIAuG42t1KzilmMVYI6etT0vjJaqbB3IHWB+xLZOzi/PnOLJrLtO0YXMaICnVQrSFKLRp8VSv
aJ+FNZBzO6o4OOxOT4+KHHOpECts9/+GLudUFhRGV6Y732J3kWLxgu9K2iM4nfret3r7eTBpRLl8
IsHrl0wXBBRmB2aMfXgbiDxgLwIr7JdZ9FB9PxsJITC9l4jWcjuLSTCGZzu5V1NikqvyhKrzZjqR
CEkbkTiO4kGDy/A6as/TEcolIkNXt/yMwzQcFa7nfmQO7YRKTFSBzfD8fH2i6z+LSiUUPigZFbSd
iekDWqqSroej8tjesTOH3YMij+Ue5acFjrmfm9/jQJiF1HDwB7F7hlZ3WRCEtWysz6s2MAA+7E5Y
k9FQxBKAJBm/KEn4/Wn7l4LdTv862rjZJnDqvrEQvo0j784NhLeVOy8rxfvoIjWRo+6OKA8n3Cc0
w9TI3NDLHQkiBW8AR9mmquARsv+SY8kxBmCJ9QQnaMF7h7vs2cq4xXL15xUa9BjXr3iGe8Pl6zJT
fjPSBCAW1Eko2VfKGVebqYjDeto/Z8z0hbRhZgeiM0lxxNhCkET/+xDCmlRZL9Ap0hDRMFF0NpP8
wzr+chvG9dBpd0JxoX/Ji619D60adSliOWZOkUCODfvRuiaG3HKQ4mt1mbNBXsgWMrRWUUWMBYH2
RKlD8X/radQGLPbnufjRRzsnT3UYBBMNAu+0JfrTqVY38EgV4uD/bdX2hxkqiXIXexLaHAnj84Do
XQhjAc64v8r4HcBk5dOPJSSQkiJDIYlPxKqC1Y+6hAlqxjlJ+xaB1phSlW7V9831nbz4wdPh1vT7
KmZdM4RwKEfr2bXTOi/ahtSLQNJFjycsHj+idCbb/+pc7Ed04bqiL69ULSFJeNd/EVMpeKK57NRt
w+zSwcZgGXRku1x5l+RISNTalDHVVbpG/uVR4GvCEn4OlzLtdRdIxR5JEMAwcTFfU8lCSDbPc9hx
44LpR2Pz4ZA8QLat6NuG76k3bqJk81XS9957MmTBRnX37JsdYeO4E1WtLwDDfy9Ae1WMLSM/092C
0Bbqnbu6ZIzREgZP2IqZhlLbvGOyrXl4bHGPOIKM6PquePyasrjvd4aEtv4h8zuKHUSwEzHdJ/Vn
zQBolUBam0Y0d3uOHjJIa6bUjAd0+7lVkkcGskUJ/sTTctrW/rE2HMzOH6PyenOTjc68zrSOOaoy
ZhhnA5s9eWF8RM8lvcgSNSlFPgr8SPqUdHiCb1CfmSIAmSJbK21Z6ffUE+ehgV7HALwdclQFjrfY
2VcqVQwgntyD/wbafuE+A+pCeesCGSSKpmu1hcbIFIZucEp88bjwFQCrT4JWtvJai3Jxf2L9Hgf2
OG5k64VVhEY7sirMBwkgucOICh+J76l8QJbgQH+j5PZ6OgxRoEfGUNiZ8sz9dR2tfRWNklZvOmR3
0NE2iRydXCc1O/IRmrQ1pdD9AstwTvdiMbAAw72F4Q09IV16HJhjKySHeBzyx0oM733iAvO4d9fU
2XimB9MFqQ7PU626CLVM6P3UW0xAsa+p/UwGWLgBJCCVs1Ny7UwKYCDHPO8aLZKFfkSJXYXsNh3E
pai0c4MnWcaSfMhCGM6FBqvU7MDo4IAe4TfFVrRcn+FpVjy9rGmlVLUh4CpOAzvjZbijX1OHY4ai
rg2TouOYG//sjD4+pKK8uGsJmIvO2B+E79YXvpSChzuSnHheiGYJNtQXZt+Srx9INyZRro1zWOMH
WwZSBmM7op/+rJKZjU+HKgfMM6RYdV0yuirN7mrEEqGTFsi8D2h9umLaX2I+mHSaHqGLVQjWFQrT
u6yepv69GdJ5xIS2a0uFciT9k+E//2IY0pvySHLmnFeF6VlwHuLqanp25B8S0N0C7HlDOp1niYOI
qvQRezjQSxaw35/uyIROLyeg07P24ZzUTBosZy9BQeXyP81Y3izb5Xd90knXY8845fd+uhJuBcEU
RIJusUUn1B7j3hRqwZlEqVOKHZ/ASevU/jkONFRnTukdNtXX/rB/HpfiQp0tZ6QQKKMlcls4+Rp0
1K1eNWGiwwLc07MoSKWTdeThmXMvGcDPK/Rt0sfGNwyMCiHFp9cq78NQ857aAKBZBINhI75Gyrs2
oxjEH2nQLXMhxDPBiItmimyDgrNOaXPU75a22JwdbpmXv00XyQaNJV6UYjygRn1Y4ia95f7NLboY
8Visse3k9pWmbLz7vWD1jShoJozZOICUFwlgAte+kIRZr+Iu4aZ322utOwLKMawCStVa9q8ybeH0
ijwpbLq9teY/hqgOtiqWp34y/+GvyLPb66nCmKVy/j0raCFWrSBDs/T7p4S7FzB2kUnQrypX1W0S
lcl53IiX5y3bXG60SXvJtYi6SDw+gGe+fKSeQ2XBYCLB7Y+ZJmV4zB3gWhlPW8nhCUc79Meo+GCk
80zpYGNVMRtLdCsI/fh7XLlZTdNQblqUi9YGeU4lwizXM4h5csvc5BVqtcQ6BwJLE5B0cIZp7uTv
A01y6Uv6vas094yTTcxtp0psaFquVmQXDYxaUPDvb0MuC/HpXViD/CDDK4XXNK4H+MWlNaM8Csez
uLaVdovp2EVms3aQlZFEuglixn7YIB2qsAvZV/ZIreitL7GCB2xiOJqJbkT35eDLI4L1W3Zd8fom
+7VWQsFA1qgDxgl+OE6LidP5OqQ9r0cf+tosZvrqUwkqbKywAYrJsRvvVzHouUqgpZdi+BrbGfFY
6PlHslYxvdb1BR9yTgN8BYBJ4puY9MW2hEgpN0ay9l1Cmm+n24sXTlPjED03XjIfcIhNvSmwmZbW
/IbLEeIxRcz/OgVzgtUtUGluOIWcHJpkPCS6zEwvG6Bf8pNVRhidizxKiasMzRCJWaxvzedoYgpC
Nou4GcoPXb5WFn0P4Kg+dw+vmIWSy6Pdi4HAoyCSpR8kLhnCNaRBu/uh1P05mcDdHOgWzPMR4X3h
+k5dVr6BrCN+iZHTChJ2BkCeV3JgFjEhqDnNkKC1/QCy9aGFfy1IFz/8iJCUUXj0aZt7KAlISmKB
/A62LKkw0KvdeD8rnhsat7IXLzW/tYeW6NPmFgk/00+WO9wcqw0DAy33yFdx3KOmL0Libfrp4tj5
xlu46guFRrKBOZ67ewtLmSayJeH8/UPMLYnllfKOO1f+GNH1Cos3RnRqmvfk2IhSemDn0vi+pSja
DIonWl2m+wVO/xUhHVDiaApV0ZcsodU5pdWQlOitWABuHTKeCHAtxI6rsq2TtOlk+1vxny9NGJEr
Q003xEP6YVuN7fINrt4O5Vb46E9Jt4RkZ9NBr7aZj+SMJYlP/LErUPw2xuZSK8nSj6DB+bKkgxtz
HrzKYJ0XLTB8Efv2RcvKGE02A2TpSUaL5zNwVTuLeQbU0q56FRUhr/Loqkb85fwtkFfaDaU7xfRl
RaQXr6Lg+vgY8VKjxnhVP+Sm/YlSg2A6kCN/SXr5v69UqpKtp2ly9ginfSaqfNqCWHfVkyjuU/U5
oCQsJJ+5BcCofs1HR3AU3qmqD8jSxJv3WHq1edZdW0H4C8MVejBlH9EU90N27TiBc9ssogAAMiL8
J382AoPnpwZkXMCkSJjZYOKGHzHFeEr/M1/mJ08H0xsv7zTJOVyOfJ8vMzglJJgDQobHdq1g9QbO
IPUud2mHiDbytPXHRf9E0OtUZjm3RDsPIEMOva1bHmx9QbGsAZbBQo8+G8vzpKW2C4QhY2Q+A1l3
e8aewSA/WpCIpkzBY8cD5Xu+zCLLTamxXx0C8TbwvNFKM1kvDDHdoC/uDZTiPWN+mltfiSB54kdv
OiGMbSTigx58aVaolV20yNa8AQMeJE460d96Xad46ofGR1n56aBXE0BfcuEut42ArBC3pB/A5kAS
JGZMBazdKTuWDJXXidUbPvzBH70J4jo5b7UBzSo0SvLPH6DkMz4pZJEEfB2vzBMQQ6sax/VFxU39
qhCqvUCXrRrblUsTwUWIWPU57nJgVyoPJjZerV6s2IAlNHd55JfZpF3g8K9IqtTNytVDTHGXCqmE
biNwLKhAA7qhsJC5VnY3EKt+DPYzQHAxVqwLdQtXos6qW6Jtmst311ItKN2Sja4IPar2Cqj9Lzy4
+E2yef0/9O3hldGdGy/B4BZlFfncM/MPAeyN4FWvdbsnxhItm+k5FpWM4z08alp38PgatMTK6Fwr
8hpculLaNbPplKPHIfpHtNhr8MiRSuVTT9fCuvwoHPaMWrXEYbL4gz9E6l+jf5N6u7NezysRCos0
v9673D5jZd2tEHNBmMM3VKogpITlcvXRd/bZDnVKXxiJ1PMJjM9jzENOxk0cFphdbdiEmhFo4vfE
XMvbpXC3vDfjGiJEmjLyGpxT/ktfmyLw0sPmfcod3Brc5RK9zORFsP9frNDnf6oGfaTzT0VAvtO3
MN2uGG32QEWiKXumTIGVXzLQIVQbiLtj/Y8gvYpfyaUlzbyx7V9Pnb9FAVg6TjBsMA9RziknHI25
JVibigK72HGSkqRJDPUOZUbcx2+7QXOD22tdShV3qEkMlt3SyLzlw8FiKG/9WNiJwAk8lvWWvO5Z
UC/LUfECqo+tCzlGnlCnjiVUb38CPKsHwwaXAi4H6GUz4KJs69LxrTWa4G1UKtt7CnWRMp+NArrr
CHlh69bxz1L4zM5SGEVp7Qcofdqqwtm1iNP6yxChnbl2e4zXefV6auGqCMtjf2Wa5+vsQvAbaumX
lQCwSdj6bgsSjaP/K55NnHe1iQ/lrCoA8oTvrRIgsPHFq7g0j3aZwHnBTDUngLU7AM99bxUgcWtJ
98wxnCGBMnuYu2kx5Bu1/7Xs9LpJTNdVdOCh7LxiJkuG0DEZB+Nwvf6euwFriNYZh20ZmU3alAdJ
9+DoOT0mSVcI99/F1kQ4Ss/91201OZ6//PYyQtOpWeh+Dt5eSQSaqpX5ICu0YbeSXRzU9ROkcsES
86/wC/eeUG1po2+p0MTzNb5tSxhIWwMNQrI7+4FrhqbcC6wqMqtjzudUymJqkJCF0yhKiGKVaFbH
xHYLLqLu268qhe7djNOOAcFSfNUWN0aMlpKq7AOkKIx1xBHcG6hgDCuBsasuqUXqjAkR2uoa3sBl
iZmeFBCmLzC2P8yXz2UC7Vc3AyPrIvMyRSw/jUC1MVfWp/ebxeDs9P4856UkdZ0lecGRSIJgiGs1
czKpHh74+xgBrFhckA8puuM0sUWNvopM4W5l0VH9XWn3m/9ZLu0GxCJnor+lufpmT2BTf5FZne0K
Xdy0CeJiOeTQP3tr+lRIqFNGOnjvJJCPO+BYvG36u5cSuaUzp6HkxHN3PaEFtumc+Z6n/r09Rzav
MQcM6nyYxwEMUqBRnwWKqLQoh0fu1W9MfYf98aJjs8Rn36W+jtP5KIJLQ8ptL+Op6CmgRVk6fd4N
5f4bQ+37IEkfmZkFcPlyTiHoJQwUz/Ojfhlxf7OnBsGWilNqzSEiLl0FKNEmpd4hmD09ImDF1qL7
rh6WoLdiKBZUS9eUoVP0eAcanmP+8eqT/FeCM7JiARBf3c/zzIc+89bogRxQ0QJJ+bYVnrlC8FIT
LVFIfv7C5JkEi+cH90kX++0PfD13PkoDO0c1WggGrfJpw56PAjwRTZyaTrNXc1HxjJsuF4XRFc1G
Pz1K1cd4ALKgV1twoUvuR64izL5/wUv4FcJ5LqDp4EGZfaThjoM6nIYtEq9dfCUi1WpOR072TY1/
feceZUoLzLq+M1C2sSUfjxNxdtiU/0/su0pASRBMkZxH5DMEY3vG39knxKt3m2LtL53NbxnpqBre
Ty3Jk5dxfegq45Mwq/5RMhqAll2w4fHt2ykDtdhre/Ajf97M7NFzlYM8Uqk8QieMA1nsJ3E7jKk4
a+Tr2m39Cix01R/iKT4/DHiivDC7FKuqZsin/VuwdCMEIxGVIe7loqGdi15P2T/Ej0IWBYxxQGlk
L7E1WoKBWnycqG5klZZXXwXGd6H1ZizGnmo6DPIY+OZ3ivwPbemh2FEMaK7glRZktWK7F8MdnQtX
scUNbM87xNhrmzedX8rgVUt2yKH71Eon4Y34SHJFqXk/OVd0J4O6FQEX2MLgurnqfrzP/Vu7Qhzx
31uxRKT2vIDpQtqbN0bFHUaVpkV/zIL/EA/hOUQbhAKSSVT+TE8gA3R8R8fWQvjZvTB7AR3poO4B
MFAQKwaqLWKOiD8r4/sJzt2SKvG8Y3afK9LWtIBMrBv995SSJJM7lTBYGsaYifKCxRdKXSxrnzaC
B6xTePnaGnLP2xqtm91VQv0i66OsIBVYQ7MTQgs2sGIcp2z3Z2I0+dlFC0BGChKn34A77Io5Xcth
7vHANjFWZO5HMvU7jBZa5stKbWiWSNvNlDcJbaNE7KW1G/FHaaxrXB4KFxLceEvQms0Y6XhobFNp
N8Wrp7iwAR2GK4N5o6lEhgW8vD6h23HJIg93DIYvL17j0E1dF/db/UeyU1LM47gbSR01q0sGBRiY
zinkxCYMkBhrKK2agGFAZQ4TiiovKP90E+oY4cvEFdOlcHucw2aqRHjfEXPpvnloz84GAF+FnVEd
JiSaLKdZDshYJgiGIiqmEGYQQqux2JrFNmjXlusx0ObRq0G3yUQZDoagaX9Z7upCbMtZZezTQ+PP
dFt0E9Wkwn1osDSx1bEiNiuMA+3zWCvWuOsaV0uGI2ZdQAt0sURONh//btsomyI1SWrq2tK5IYKB
e/KaRS+M+iI5ux/FCMVd5A09ZI0xF9VzwqTTGq+80FiiBcTw1Nnc1zAzPoRMx1rbrMnazX3vCAIi
VE/yOnJ2fydMvCj15IO6pQWzQ4cwHiriIdgPTzrc3jTOAEK0NLMPMAP9gHYROahHn8MvN6xI2W6x
zd6ZfB17gzWK1jKC2Sc08761F9CaSegA/5fRxGA2cQj48BAW3BeOITaE4J/jBi5q6WREyAq+Whzn
HlagF6arhJDBZcNss5kPmd8g3bzI0L5yRLlSM/YyrmOXpuYhAGlslCV6z5qA9bWKkiiYNEAduEOr
zdPJxIwxVZAdu6N9vuURRr5LXI7Zg/FOPyDczykSmfDmIeVUn868NMGe7lcHSTLfdeNhFyp7uFZy
RWUgYQaxkpnECCGo8rxvj50vWEinoOn5tWivJaVbBZ65NBquJTKaKIrZViiM5nOPMAYCsXZzVpmp
FREO4geLvwmWCyvdNSFqxcMeNAB6nnjAlmif/+0dzoBELWs3QLRR//gI2oy1+dUAUlTtS3fxxBK3
HKhC+YP15MwsZQjBx0ijfg3eWzfL5Xl/+aN9Wtqha2pqsqpzS7SkbfFDQaiaI8MM9eahZ7WC/jAr
S3tw3RAC8BGqwjb4WGkT223+5AQxuNjXD3SAw4NqWUp20DqXfvldF0rhmSSC0djjTMFZyD04AzqH
nSAaTu6bOb3uIXnhAxBHkCzmHRnRqJlNu4CK5ZN63ASb2uFGdUgH15YEVKUfEq6YraL14jOiZfAl
RtqEHZk0LhzeqG5tQ4VAYVVaiT5ldeS49Exz7bwJZcn/FXFIoj7BwOXg3OyGODy3eVrb6bqwY09l
3AQBUQKIejFfXGF/YhaTciCCqvt4P2EN3hW3BXZgvF4hqmgksl45s+/jC8mWpUSk4WwGjxFEc2gu
bglvHaAVSFNw6FP7eNXX1iI3+fmWM10k31yevnEWvIFYWHCcH4zTkJlYtYBHz2gPbO8q09aCakh7
o5R6zn85HDmZmUxRg5qdCRePkQsvJAvgVSjrT811DQifAi57ru9Ufb0hEvV/e1/PFmGVzMIh/4cs
SZXOGQLVZwIyWfmq4L1OBnbNLKZCvz6V0QmOSSXaFSz4UZ8tiv3HPahNEWLmm5xfqAzYedHM7Ykx
65QXTOjtatsYB+Vp+RRiuAGzE6Lvscm9CETLpRP5rFBzGSbXGTqrfB37DdTgpYOvNSWNk2XSS1RT
+AH5yBvq4mCUZBEv58p7c5lBd7Bibyn7NDXcDJP2iDXL8Roe4Oa1s4DCPXnIjCmrVVKTPkAwg7Je
0gQaOJVkj/8mqmWRv98zdBNmirBhRoR4s+p+LgSLaV8migj2hyxM+9EYU3QWXxC+Va/fGPNntJ1/
GxJD/wbwqQPoa1QWcheKqkd0j37StlKQK0oBL1YJSAcZ0vyInG/ikRs1Pdh0xDPIQzkseQ9JC6gP
m58Vf3jnYGKfVOsS7iHPZv4BrVFJSZOGZ5ehm4FA1s9FLYWDKjJDG6hCgteRXsnIpuNmKydkUge/
i75pbxdQ2cu7mLVkOCTRpU5JeyxmAzsbRLQCAlxc332ImYvbN6Eb52s8+WBytrJDJB6Q1ZBzrpW+
DK9y8WpL4XoQeAj3MhnDM2RKWIocr3DJSrWnTB0WDORd4YMz8j8ebsdc7c3Q/lLjdeByAP96tx6z
myAn6L3R/YePKo3VrNfg+OEcvfks66DqbWN4L9lalS9MXgey7FbSfjq4oObMGWk3bcoREOr8aRpM
S+y6zy6vwQHBTHu7JN8bXhev2bG2irVp8pOrCJQlgkDPKdCEaPM+vFviyKg3g5IQDR0BLzElTaW/
ham1BEsSWDYNwEsbS803Hv6g6NAxrG8YOZPfi/mzkk3HeYjEbswMdxsMeXiKUSk1OmaW9oTP2cjZ
n2hg2z9w2GSoMaWWn1XI6hqsS+TfZqClHgX/L9pZhaMVh9cHciuNlDNIarzb9wi0dFFP9X3371gD
2Gfe2Tx8NFQMRHriafatpnkW5HFcjLOLtgi9EHfDyXaR4FAqhS/HKwBeY/SgVN6pRZHUc+iO9lPN
Myqjctsfi+pSP8cZDNmE4X6AGLXD9Rk1lYMquehFAjnjxGCzCmokZ9U4qLfb7ORFfbEgKpcN0bDa
eZGfOJ/QLMDYlVwvqATyJ2eebubMacc9I8bR6bU8lFO/AbxbvqN6E6ZigyD2IulSqQq7jUR55wo6
ciL+9Zeja4I1ZnjS+gPQTaCCNlkX/MWHNc+UCZU34HCg9w/TF4MgmprDTcHbNE+IYA4f8Vmve4ze
2Cgd7Ic0qnTd9duZxMLGqgFChEVn6sNwZbWSIEwrdAF4nYOPOsu6qFLnpSrb8HvhixMOpZ21yXRS
Sgs2ZtEojOSo8rG9t55w5LFe2KzgHT7OqEkFYiTeBbGUMVDkIHbEKVSDgLAxoTvH6S4sjha2BN30
ctYjVpeorxxP4rrvU7WvVBTZ2zRbS+tGjQ93PJm7xM5skZIlf0KK6rkhcLQFFazIxOfUVp9qJzD5
V/iBPyPfsT5PbOE9ZRgA/k1wu1jSeiIKws2QUAeFdbEky3hBL4iB06+6mgdoDkBwu2PHhm6lRgVJ
n+ZNaBSqSwK/9hYVpk33qKlgYIp7Jy+3tmzc8UGD7nx6xLnzAtqGBTe5qqq+xVuCArbhJksFCqHF
0p9luClpT6zF47nf+Qh/gnGn/bGc9ysLK1hZRj3BPf9O7eutaOb4PHoVP/0o1y+3Yfqo+H6eWA11
LteTr8Dywc8NAkzZI67mlU3Wm/gfysfY8OovYUK/nEP5067BEHOvpMwYw+4lpvkQ7WINsy0IflIn
WzFiJuioXd97mu6s5w+jPSVmpZhsXtgteP+eLPsBp8Y53A3+zpFq7l+ITt4kJFJqoMiFX8TlOzti
vgfUyCb+wxD959RU2lBeY/3LDebgpGPsD48o+pyzW6oedQywfdJYdFivN5gj1OFqh/2O53uhr9no
1h51T9DdSuu/i6gSw5wTtKalid2rZCVQVf1QcdBvqpbxJHIz9fxL673URzrGfj86dOwIlEDAGUC6
+lgkVjbmvsZOfEXgwobXGdVOh9DqLFupkKawINUHZe1Y5VVoWAhPT9mlZwp+uVS2Aqt/6d+BSizr
4+10/HqrVBq5LkYgwgESpO3byehMFOeWzay+d06bUrdrBDwIPakFy/pZOQqgPt8U/ucRwy/0cCVU
fumunNbJTqhkbJ8e0JVr44NftJuOHHQPMDh7lF5hjtR60ldf+VmKAzMUSn4lAxQxzgZB8QuYIFXT
iGnUfhpRKwtptQUF8TO6HUxLLaYReorrlBr3nXYyhdHTZvCIHsYWnz37QdZefIio6xJ7cJdapHV2
Hcpw9ayGRxLHMCEnDz3NfGOF8bSACXykpFPNQiucFYGVWzUjfvJ7NlMgScwfI49LzWWKrFBM2bo9
0WgH0gvHnvLzrwdc3hErlRL6acLp80/T9AlkI3RLbYIOP6eLAxd6Z1cVyEPHwdLFA/8IA/99dueN
dSJpIg/MzIqSGVAU7WJcMhTLquUtuJGzUs5Zcqvoh/ebPT5txKDDdcN2myw0ux04b7JOfdipp8te
kr9ORjbH7DcRYDA4undzbNLU0QlFHMWztsXIu+0QV8M7hREJE/IHMGxB7ZPTpr4x90uw5YAbj+g+
YGspzHm+tsVexlu+tFrDFNdpUhOzs0Z/j0wZ25U6zrLLgL5VMzogaKEQcV/NW1QUAjm4j40SqVR+
dt2eR+SrrCIql/u4Vbl7CLGsW6w0OHDG78bQ3eLTHRvAbzvAlCIo94BeiasVU4U9pnOOp7CkASnd
iUj+tu33gvnBPos49MYm90Ykur572eJBuf+SZTfp3imofDkOrijBTyoi+K0WNCIFks5Ci0JfiERO
WheCp2xj2yOJ67zcmOt3ujZWmQxeaWaggeXBfgARbeg0fZuLwe80DYfzeo8nlKKdxex22jtQNOLj
IxiRWY/3F4Q4F2jV7m78D6JcNNwPhJVWiCoWR6SpiyAnk1elGhhTFhEoSQ/XqPqcZP6Sd1h1qy2p
RRIPS4pj5JFdbqNhyXU2fkTWXcBl1DRbM9dki80x9FiTqsE+Bc0UJkJpEx4ufTmm5maaegN/g9FV
B0zFKXG26us7mYFo9LCwNKUO3nesiZJj3KAGDDU2uLSunN5raUrsr0mMGBKQJbgeIY57EBZUuDDP
Oo49EzVNAgDMViAzF/W1Zq23ITzcwvxbCbvw+fRD7fikA1Qg8oEe/x9pKOYchqkZ5nslHnYhtaoA
ZIVNAjSs2cFEAZoaUmlv8DDudKL7myZzK0ATO+8gj4/7D5iJ6vilG5C3wkT9ZnD6JNbUUOP4xq6W
L/Tb+qJ/Onr3DLd+QlIRFzlRyrgaW/zoqm1g4mXgBvggJZci4M2yF3hPZL3/pm0965gXwcTMfLah
Rb84L+jHaKsgQiogPBpL6LOc3ts1AtVa8WWakdGjWuhW7y0weK9vlsShfny08mpZgp/HRxZdQh5l
uOFT4WvBBrcsZXtN2E5x2eYPq1SvxrA3umHQREpgFCYF/swOsddnLLfB+QM+uc/vZTP0wUZhb0BL
BwN/u6oRNwcxK2WYXQymZ24s33+WhbUu03W9ymbRG97HCxqmUbYfOI9NHmnuSAIMbgnGnHTxNIkC
9azDFLytflqfUDg2m+TbTo1eq0R1dHXYT+YogEan0hRGX4EJ3Sz6pQHTjZAZWCNUYj2L+q/IEFg1
kfxJXlOroYIFKIi5JkipV/UtgZEvzbWjxnCJT+PAr8sWVoe3hK6ex1S8TsE1DmzuzFUyvNyXSRvx
/ZmtcBjGxpuajDeo1TcspJvE8jsOK7Fm8zczP9ECg5u9ToSprqwo9OH1qSUpy2LkwCcRbbKfYLVh
rVab6HmJekOobZyJ2EpJh3a0gRIhEFfsRE/1LiE769HW/UfCdcTPOHXBfZZ/qxb9kQTg8OiXDbRp
h7lY8QCtBs+RPopqQxAVDOuXTP/qmi85UdMGG7v9j8NAsT8ZBNrDGv6lBNJpx3h0Su7nS9jhNr2C
3koCtaZNSvvjS0UXPt03OyCPxP3nSmCS0qvpjvodKcs5/r/C7kPW0Ez9dny/npqz+/asZ0XAJB65
0hNLwE8rwMV4Xmxkhs4H54JkXbcnkunkffhZF5gzNvPzEtVr8SNfmki+yKsYnjov7yUHOvraTeLG
VrMerqOPVzRB8iij5zno45nyFBRKSiyto3mBv6aye1dVkJdc9jG5a8NrUfyBNxGcNZrC3qmqR5mz
fbQXBuoqw9quigHRj15V56QNSlBNV4wo2Po0kmRTR+yq3UfyZ4nJRb83V3JtZjOhcL+N+Oi2A7vc
q9diHXr7y3EYcsdMAdTJVITwsxei+rz7dIWnR9IhAc8fhJG/Q7v/OK6ZTfy/z0sXN+z7pAxmYwvj
TckUrqs79vi51+ZuFByA3sHx7ibI93DseN+cVljusGSCMvdr9jQmxBWdceVp+IQEglWwUGHaVKpR
ABXxyfx8WyTtDQCLnw4/woAxpaYi3WTElGoPGpO6Y1FYWjpdbNJ3fQ/OuRa7wY5QAAJUZ2U21U4T
plhDXDVGa+ibW+VMEZq+CzptyNJzzG4wE3daFavNBS2ALTjCens+KIw2zboDGwRt1fNbc9OxPwCI
Ujn3N9lgGlrO9+DFWpatXDyfw4uMUDdwEBOZO4C//3xhMF0gZNtKCqgLF5i8P47MdvWKf3IS7AkA
jYZs8fBgDaLHponbCmZz7MKPIN6SbIHCAyUzuw4FmmvY/NPuVtzVFqfuZOXHyLhjxwBB/PfV2oXA
mJbkRkUoiLqLIphWAtph1O8g1VJyEPg0eWRQ5TyyoH8/anC/rScx1tFAHDxT4VHUyWSjINUF9vPH
j66w4PyW/lIbzS9xG+vXoztrHk29kKqSIUEMcpmgb0I1MERVNPeRoO9VqL8wNTRRYKg5+Fcr3zUd
hO1pP80+bi4NpYfpEhsdmzskmGoOnsizKqSauY12ZHYekpumiMuvHCKvKcxdjXU5aD7M7Dm/2nKy
Ahh08g8+CI5ojDGjhXlAfiwGQhU8JiR3AS+lAMZBS1/c7GbQHfL+VK5SYMbVhedUv+FPBNvDlt9Z
EObzhUj0/7x97Xs1cA34892M7VWZQiPv+91vsd/raBFT500byCkwG3x9yXpD/f+0la419V8Za5ws
yVYRFO90E7QLSvIuAjd4YTnjBG/h1+grz7fK9YYOvMtwR9EeJceDdk6MsFckVYr8Plvmo4MHB1d/
/dqFzm6fl9nUd+noUKZ7XEUI55fTd0w8cZ8W27xpqR41ntLvza8Qrc7RnrmCcKYzr0GSSkYGpe/W
cZF0doHCzdQ8WgSOmkNg0614uFxsUTAVp8JvciiRvOu8yyf1CVT3YFxzT0CITQgeyzs4j7WRPT6o
4sYMQ9KEC7T5SVZ8bySag4jY6jhUdlyM6NgFk5X1Lypg9ME4RiBiEoWQf3R5OYQDeQkciBE3mR5X
4xJvu9xzukU1zftjb2vv41Yc/mS3RUqXl1DT2k1GrQDDwnKpP1Hrh0Dtd4mHedr9PaQusOLqoYE+
s7rYmR7BE/pM+c71GwfJMkQfWiz5uFwoFTuLPhp8TYU8YvbW8cFvQScSHz+bcXQhQYfeBUgU1ooX
jrPpMkQgq4e+b3kd8E+6vJHI0ak2ARp+x0q5l2ovis0IHdTH4OiBNq98G25V+Rk9znmU9C1jYuBg
rMlFSjDVhXhb0EX2sYME6qlYs8MkkyOUlU9klIRR2cb5fhvZnUJXfFvBm+EJOpCDNMTfbCHb8RAH
i75nXC9+rA8Kn9Q0r+xW/e3Iu3an0XzXntHQ3jQHjp1IDv4if31khG3F5JxW/PAAfZis95M2GkVF
HNUzISUpH4kDwYi3/SNIwYp3jHK/90bSaBvNfTR+KZaKe3TvHlrwm36B77yJAgWAsk0bD3iw4Xc9
UfmONzXudP0MDxZg23Ayv+LqfG6nubRUZp8FC1D4Jt5obgLLyjGzfr2Z5XbDOq0M7nZOznxZWY++
piaEbKtTCKI/542Rch0Wrs7d9WxzCQ3MvEzjRdagEsqf/CIrnJp2pWnsaCt1bqVYR3a00VXeFeEM
RTGQ4LmNS3HrfS55etPmMhOgaTVESMu5WM9sCLXzDD3SuxSrnydxbYFelwHqqVVc6U8KeNECcFYb
rB6wtRmYUqyQDIOuQn+zG9/fzoSEs3DEtlw9kLsCgF99FKq/ZQF43y7FysQxMBmqrMNo3i67Ujx3
KO/jk4TZcVTvq79kAyTbb5yttze0eq/svXMzYxzI4PnEAy5Sw1Dvhj7EyHH3PnOPgt50UkXzoPjc
8fLzzEkSqsksAMNMr3V8ODB2ItKp0EDqzndi/hHAP2EFpEaM2KSVwnsnJAmYlzhvpKC3Ryy+L0kD
Uy4AUB4ayMVbCy4/Uxmgug1m3KrFlRHjN2haTjtjCTfdr7GLqd6hxHPDj1TwzIwgSfe2iGIrOYOs
kHOzzpDJ5kXK6yv8dvv6P2ysDareBK7EiflQ+lqX5W30OTjpE1O8CAwrlN1+KokyUOFdWxe/0OiR
2kTwplLQ9NtiL4cKnvQ9sB+aD7MoUfHqyZOwMY4kBT0CxnshWnbWwp+5Ri/99r7RcyypEo48KxDJ
4IUft/EcKq5ywfgZa6EkzpwbcjS5AaAERz5y5QBUzvEFug9iTivMWlXF2yU1djcVIB9T+lf70kZ8
cpA2ch0lUjHNfyoke4QGbl2mhP1Sx4v5jkoXaUZcjWSjZSUjVTp2r/TEodnhxARE9FmIDuwE/7Dw
odln2fl3wlTDEO73dJGFaZDvA8IcZiOCcyogr4Q0BWlhpRMulL7QI3LkqjAQV0YvCZYHXCdDoUCp
CjCvlThKm3nJn9NudwYFl66jbMUcgfkTkcxzqRIH9DNqCyS80HrjTCB0lYuOOz3iSwWDGJYEY9xe
OvwGQ+8Lb1e4zwlVMmHrE7UObUtYyjjWYKUcz4vjC5PuEFfLXqTIpTxmBlyL8Lwgfd2TcilGTISA
P3EeG/0sD2M4JDedrytvepXSCkgotOvfrp01La1MeU56nRuQPYFmpaFw3QIVQh9z3Wl53OOqfyMV
ZiTU/J+Ll1uvtTmYCvJliymknM93rnZy+G6r/gyrrLW9C4ebyhmJTRQVpl+S7Vo0Bg1xY//yAN/k
Vj9bkw2BYRxTUi5r1xyqCrwma4QE5cAoXJdL4u80rwhvrOcZ5IB1FcMHIWzq/eEKOChZyTd9XaeJ
jbgkfiHvrwXpOouUqX+Ixzed7iz0nj1xYeW+S9hNRIpJxEkaZFuvlpXrXf2AxYahswSPTT8nWwnw
8RrxhispqM2A37QzEZ0Xrz8umHPXRMlWqycU9sy11feyKrw292cotDT2GwiDwcPfUICH4LOahy2+
1iuwqaNUkpKFzfc6Th/HYL50mZnHzvU5FAYEp6fwKdVAjEk91OgemiSGyIV69Tkd41TQmj9Dj4FJ
6yz8jpZih7A4p0D3IBWS6ypdhKQjPnyrXaXPQKYh3c1GgSumMv8qzCD9LXNJF/yNDXueJEgp4Kdn
md4Hx0vJwaqOSw4Y+RyuBEvA7EyOnZ0WsAcKAMbh8T8n2QjVK5Z/JLYz4Flnpag5MYzqciSBvTmA
I02hlu3HsFpTv7ejYmC+xPl2uAGDf/p9TvMZNWNN6e80IzSyONsOi9XhlUeYSqZi+fZwdNVlL2Wn
3LCWI7NvMkXYKxyTGCvYhUGbI2gV5mLi0MbqSPxj6tgBukstAtsJvPzrljfwfc2qrgedyTVdX8S0
7NeygflTRwEhQcrYE3xcu2/87O6EHLw+k2uXeHFSnjuVFYdgj6iId6PDlT3CDhNgLsz0s6H/1ShR
mZqy1SCyT1q/YdSrAkI3IPragKdy75giqa1o5bBQl5jfAVbC8SILC2csIyzkF5a4MHdYJFPS5h9z
5gf7UPA7eNgclAzaGkdBAEmz01PHyGFwdw2YEV0x2GHR0bxM5vFJ1Qu7Cv+0iHXBs3MhEikTYooe
ZmCPKB4ANgcYWXUwDrAIWLVSsPVtN53LRusLyPkhVYesGt/hzWfigIcIrQtWGIOjKY1v4aub/Er/
FF10YRyQS0WMSYd7OfkfAPZMzuZwKEnTUA/aN9NCRr1SJk1BYTA8fOG4Twtok4V7sHVc7KGRAqPJ
deIUj1CnpuClt+qIP7KJyabrZgoF5wai1Cf2T/CUCcPgon09nfAZ9NR55nC4yLXldggnZ0yQIq5K
etKtKjS2av07QePGx7QovCO8LEarye+YD3zlsfRg/JjJnUc26Dkb+OFhtdUW8olsvcNVoe6EwPfC
33E4QEQV+eJJnraCP7RPekZcZaQ1X2azFez7QBsABKkN43qpUhdxgSUu5xWgyUaK1QGgTsgEEzy+
NPEGsGh6A+5fFLjyeQOQTr9W+MEuny7lwgg8EiK4qL54qcDtYY1gPc8OtKPE4/MCqzCnL8mh2M4b
QXEp9YsUmqMflpsQ3m7MEgfJ/lzgvOZ6CvoxQJzezzL32UDDr3VtPjVoeEz/CnKPNV41OscddHUI
t8jlkEebPn5iOqaoo/Odpjt/24hA9xoxmmGVEu1lFK349kmXQXe8/Kk/cGGsMVFNJSZpebA8p4o3
2/p7+aHKRwF1yu9esylp63h0FeUEiNmP5d/GtNCtBhYYox+gGTlnLZbdZopXwjPIPuiAcHoS0tzx
oYLLCKHk35wMLBWftnI5kuGrlVOupMcL20qwO5sFJl3g/zExcgkYrtqSajdDzhQ+nIMZj043IOqU
oYA6jBqwP8UggL6ZTii2zZZq+ACbhXIRJzuQs42nSyQXEPWidAMcsbsNt2L6+wg6ouScTQWMZE9R
StKDNqOowuj8BobtPm9G7D9H8kvuxBdmzc/BxAX6YYlm29y2Zi4iYfJdSEn1pyBR7wJB5Bb32mb/
fTO9epItVSx7K0MZk1/34pX6zTtWMoLScXZ0ws+0p+HyjwwLfPX9R22ZL+D/kypETgF9/bdSDE5c
bWWMXoJkPDPpNr6T2ZfIwwSdCDhAEZw4cClTsAarrsJQ94+ygQ5I8B9ATvdOwU00dtW4c49Zx8Ka
iC8XEvNUOHYIBPtQIsASrXGcrMUYq000Oqs147zADCp9/qV93Yo/sJMx3tBbbUsY8qLBwy7RPJlo
1uXNxs+Lg4Am85/qMOIAG3QSh+FQ77QcPpAK4oG4CXJ+E9sB2XWjZ7NMHMViF2/HhP0ISoW2TKta
a5xMZmSFtl9ePusDlPihltJbEqS4XxYvSjQv70rHil8VeMliYKRJ4AUdAzwYm3Vbn9UmIkLMW+BN
2xHk5t1oYKLNFrPM1QIKxemEY+lTC3ZCcq8KsA+zAG35kB/kYhhSfdzot8UHid3PJceSoXrsThVo
pMersTvrclyR3T0OZBeXblkPs7PkWhf9X0A2C+c3iIDoA90uExLQwsJXnb/r/uDuFyvZqi+Lvsoc
LVTV5Cx3V/h5kW2rpDV5cpKV3BhlJkI6r7W9Ae6eXR0Q3DhlUE0mI2b8MxgtoTtz4uly4aO074vA
xDWlYQPA3yUJILPoOL7qWfrwBXxgEmp5JET2p9hZ4849Qref7smbcdl3Mw9Uw15nmxZat4AjOWqk
mL26MIytsEKaucy0JW1Fu+PVkFh1aU/KjLKkzzUZqT5WSaEdwD5zKkch0WrYjL02Ezoj6gor1+8a
V0WZQe0LWhh80w/ZRUCjgph6DzPpm5suXCGj/EoOc5lH+Se1KPwRWtcCoBuFifZg8Oans4fDbWBy
gRvd77YoIfADC9sdPJGdUiIEsmUe5wjzJHT2tBrp+JnsDyXhtbX0fpXB1Mv+gNiETvYbJQVP4uFv
/8Yl/KP1huk6ghgp6Ehz355wYbLHOMQXc6ZRYMs1q+T9CTgOzixbk0ep+T9iHVkSqrBsrvsxT0jA
J22uIWsv5zSl31gH24TBUmkeI4D5BHpxEOl26187WpfiQonMJXY81tE7HnF3/Std3vf4RUDBMXje
537kszaOcqoYZVZn/QXTpReJU/StQpxjQK8fpxTe3MWs/a4FYqCbvkX8Wl025KoniTlIcfskpHvD
mVoQUqZcRmeNSB+yuLbgW7rDSVartDpsxY2Q0s1Bx31OWSSclt+Kn3Nn8d8r7k0DrVQooJ3BpP2Z
swyjnN8S2m1vA/MH9xp7x0ypsO4bNJusZvwHv/dSaw99JcDH9ORmsol6Q2FjmnfueFOrVpC0mJag
c9NKWpSMXgcCn0PRgmkG+Jiy8GIePl72xaVFJyeTHjnSyYC5biI1hwKNAe4oF+NaH2gJElCo2BOh
+0GmG7DWz2myKyCqPy+k1QI+FuuzwQLQkNR7zZcL97t+lWshJKDIhFSh3o2Qmxk1fq4mUc6hCd9b
jkBL4DTWgWS30z/67QBFuywaXOldravghCibmYRaU81PlHJHu9o7Lk7KGhU1pH8RibimZXd+VXkT
q0rUcSiso7xZyDNCe2+NW1YA4ljXpBhtcIweWu0bQyu52iviZEhNHv/rjqSNSVdrRSH01n6uIzly
/zyDC4fRZhYrtQOGOQjhI/uI+LU1hDEiuJFNH64xNQGrWGa6uGuTXaeh52DDIwAztOeg8JWJWrDH
QsYY8q8KzYvNCPJlz5HjCg2HtQz3Ygj6pXGjhlUy19GnzhfSHD2TTHGcY2Wj0S0joZAxKFGd6BDp
DxsqsGYkjvJRsXHA/dveI4UzlnxeyZvbpyxxnD6Rj8ObRqUW0k8PMojju5mbSMzH9H3sQudIoPCw
HziFEJvwHAoO4010wlRoaAY9GXPM/iWLb7I8gqmKbmy+2y6IyK/Ba9ohypR0wGSp+3Ht5E2UXaI4
csVgpgbPTUFP8zAWnBUP82otLDukGfr94ngtlgTnVbeO6eMzpnzGpuiOcgCclED6oIp7ldEHAq/C
5maf80dUelP1F62zNJPcCwHGP7WHf9CrJQyNFj7pKgJOJeyqii5BLUO7JnOKCaj1xsITea2ZFxg4
8c29EKcjMxz6pPUHs1A1Y0GzHXjVhUQrYj5dUSomlgAkqWD3HHEmpj8fdZ1tUQumIrq3sNVQYp+g
sR9BkesCGaJIdJmIFTZ5DZG5cbQhs8DzXRlXtjwwXaFPABald0uaz0vAY5qrI9o1kW8PK779w2VC
U3xb20llxoY8e8klT4OHmTtuFkOd3r6TVLkwUFJ/wrNIdxlJmUkZCw+PNQH6OfSBijzK+9td/7Li
9KjfPr+yXZtXZC6/emQg8SbWisNIYwunriQzkAyhgHVuWG5w4j8j+T1xeIMMqy4+15WXf+GF8wXc
SnUh7C89LaM8CinTlvZXJPot1yLoKwZPcofXefpzJImMnlkzalfElw9XMNixcPDVl1cHMXYM5/xk
Sj7PlSrT8xF5Vda1x6JygEy6G6HdpRDTzcP76jzvGB6j2jHK9f6hlsVAISqQcKYUWLirg1bjQ0bm
hW8qXpmnzV8HYKfsnb+4+AuxkI4z8eOzd3Clk8iBUh4tqVYRlRKDUF4k6nzSGbZECN52oihERTXJ
+eVenqXqsj5kBXJcJ/q2y15Zl0b6eQB4aJ5pbYu/C8kXSpXsvOPEFLK77Kq8LNT8YczcYDU5bt9f
ZPkhIO91xBB05hc1zyxLyp5ZwBFWWgrkbVrfVxfgWomUNHB2XSgccdPd3Y6Mz3M6DISQrpWphHeq
FzND2PSMWNynO/XC16h2ugtAV2SH+CZBG6aFn6PXET6pefWguLnKOyOpX5MH/q8vAsRs5RP7uFMq
cHYW/zD/tgsOMrXdm/DsTvfea3ytfjgTmy2VxE36SgfH6RJXq0sxkMNDenT9fcni69fUQw7IAxuf
NaHC7XleJJI++UhhTw4I8mZxjvN6lFKi6bZN17xJUFiMjoIGkp8Iqzw7bGuRPLPY2rucMKhES6u4
IMBo77S7Nrqb/Ib5Xgl8nCWkmOtdA1GbCSZYt8kZm5IE5zuwjDF1DW+qvUkcGvTybx6A6LB9sRKL
JZvOzuwWFV/+W9wZKquTicMsx0Bt5TmCm13cNSET7Je9KtlRuAAAHJbRdUT1UFLf3Eg938qnP7g5
h8sWh8LOPorrKYwobOQdDfF9rEWhGzXATmERTxOmr5Oe4rDuEwXhklxnN0i6Kp5BW4YDiXhv6vWv
f9racRj7zktzm7tSHw8lyK2H56JQ+aeGZuWIyRwofv0jTpr4CDJPuJ62KDziU43K/cKkmXCqRWy7
DEVqkkoq669ggCS+NUPtU9OnKeYwELl/aGTdSF1dalchI13LAeGb9xmR/ZzfNcRKDyuYXzC3hVID
23frzFry5JzAdtzu1TyzfK14j7SGc03hLVBLndH0cRC6IBTwnDD8MweV0BOez4IYBoPOffLn63GB
6uB7QjNwZY0reoeB3yjp2yVGoexdsUWE9hUk7ylC53g+Z8TletVzs2+8Ps1vxO/YPmDTdNmEskM2
gRrpUscNlcVS9JvM5QvjW0T+GRmNYdin20VekerosS0bDOKBFn9SwIF3kKoPLLXadThTLTXA8Ozq
QEv0UJLGn1zv8ijp5WmlIVWflqXf9EQHCiZ6mRtwW/ovPygbFy1FLV1U0DM4Xy0EPCPAYonc5xYO
Sm9qhoFhLw36xzFLiCVJRHrNVW68BEzreD5QD8GfQB8kAoXaaORZZGmhoUA3ICuqjHkHj3kMWgTs
c5dpXZemCdsSrsqfhN5gS12YHNJxbaPkoC12ySZqwG0/fg1Ir3FD/wAyMw2Mwnf4NsHM7p9LUX9j
YnZSrCDsZCQmnQgTAaztUngWEgOItkBl2sQWL/bowZ+LFv/ui/ka0shmcrq9YYifm4l1k6X2k7o2
O7jPiN0dc+bqm970zBlJpm95OA2BK8ZyEjf7LtVz5qkmqT54XcoR19Kom3MRzCSr+iEzSXYzgnMv
llauH4gucrmZJE6fifu5uZCsSdKhYbHL+jEPd6a3V3Hu4GF2ogXw0xUOb1J/Z/Ff8riuO9Kc6E5U
xDSw8rAKkWMqPKywfTotTzGj5PU9i2XLM7oN6WJhW3RESe7FvY2kj5gSR4m5otsTqOdMvKs6ApmT
FZGWscnUW/7Vsv/8dtHG9HX9jAD+2mm5J5iDQgG87I1wlaeD8l9xjlFsGDUFVfPRlc/1YA57Iq+w
fwu2wS9QMWH5wvNO4rQ24CUMlahzGpTSALy+aKVoaeGulP18bCIRUkD6KRg9G9dUKhLPKreryVtA
CSZxn9QaCLKLahIe1caPw2ixH061BgghTyVS2U8O2hjLDxcOAmOuUIy8k6NFePEpxTU7krVBHLEf
Xpc6l7RnMuSNkk3KoPz+LzU4/Mu58D6N9NcZiqf29LQkqs4A6sBa1DnFCUBHv8i+vtRfQgdexCbB
a0scw42BtOumxNNZq9Kht3dL1jpA/JFcl3I+sBxTXg5f9Sc9ZO2QGOjQ4FYUAVSgPXcHuHWXlyxN
HYQDGle2AHZaUyiBV6iLRpUGWLca69JGUSuMaDS2I1BNUmTCI023XeIXpHFkCiC1HxjkV320HURq
//IKPsS3E/2iJbGwbr38ZfDfPGAbsgveO9r4nJVnd+e8q5DOKrjEVCpQ4uYKrzlTeU9X8mOTAkhr
joAcXvNDvs/gBjmgy5Q092OYbqAJBWd7LlIpG+fc+yOymfBzhHrqGLAwsgY/lG6R/4u4yf4n7rKj
y3m+Jad2hv1H0jEncK2E9HUNOk3ggwdWsmsiDAPpOxnr+IwpFQ5SOdL4RYG922HVLWzMzHVK9Lcn
Xc5qdz5FqhejAHkma16Cd0qG8gVBNcdQybdc8d/LJRLe7DGadn63I2ZRrig/RoLk7xdCZn+Us8S2
/IwiBvJHvf5wg9QZ99MQooqsphqpK1VwJa8h6iO0rlSqEkxB0nHYiRJWITfBupsK9FyLlRKUAZBo
6r4sxA4WIrx74JKz/6DnyxptAF+rR97v4iLZmWPOffJl/IJXWi6s+6OEhPthtGnUgI4irmki+5oy
9B9yKCVM6KCD0bsyDIOucN/DDWAqrXFn3TCN+z2Le/EsOeFbTdGhN4VeFOU83K/wr6BV343AJPys
Slfitz38dcYKaHIXFieph19F8+DZAL9XVWWi/orr3XoxZV/xiVPl4RVXjxZY+HyN2YmKSziKS+fa
Ozlf96EVFQFg4tGPEFEHCo3n6AX0QiwcH6ji02gSfnTUl1tlzyHRIGst4nT0snT/6HSkabZKmSOy
iugPSPURMbPcFlLVSsVRuhvcZor+UtNSsfesUhTRTQOi/QpL5cpkEjUZEjfBV1E/0pCAZHwIGe9F
4ZrdZUO7PVNzX5T61uNem9AxA3//dSzN2RqiaxmyL74zS/COii4j/k+hHYvSaNvtF9nHvG5bCzur
D5D0/guWoRogA2KN82Nmczq9ljbAIHm4tK6o2QcXlWonvS8L2TiqLXVwPKrwa6u/lB/yPXExafwS
9WgvFeXXAEG0lYSFXxI1EV/6PAWB0MCZ85+NPHWpqFXOMkaPdrDJKcFebbMLaoJNdGoP3pVu1LOk
c7ERTiDY2LS3OvOpXSWtS+OXXNcrR2tJj2qRaP26YzuyjDi2DwY9ToTGrARwIcIlUhWcQKIFmuuB
sskO6HMIE+IQCmjpTq0MDzQX5W0q2AfIhtxH/Skm8K/OKrrIOpXyqNwxR4LjvXeId9kKNpFEmXgX
SiPAi+4Y48pbXkX1EDITP0zVtTNDcGqHycG5oRcLAs9kS7NlEmJBkxFksb39fGHuiEHG7MveaYRd
kz+0kWE5HtPJxTOO3bp1CbB8FVJYEGap3DR2fgInHN6J2avJKZyorNO1LONqDN9Bk1buZtbH43Me
nbo0YpSd72vBjzoJgvSRhW0s8gNbyKhc3jp0iMmJmBfnJ8t32nkJAmwvaN4usxyTl9JAwRXjdgBN
LlrL99CgBKjb0qU/GOU9+h4C20ZxJeXTGFdn9gcstzryXzFrEwFf7Hw9cJ126RrLAdrDgP0rjIbT
MX5spvdzz75VPw1d0PYvIeyB/+0/69EGcA0BFGVQ4n/2UBAteICOr+rCiDRtd0+aAkMDtbM2Y9ur
pArifhcfi9NO0QrgMGhYc/1JtcGXVgxaiDUokWyJ4VHPHbhKgzCGvAV+QzDClRurN2GXr9D0vL+V
2+laNobQj7OMAMypYobWw36e/KPu4O9JU7TUDi8KiGjSXL7/LzkTdW/tq7VcDRNUeaNpiERM/NZQ
fDgrW7B6FCVvmhWO8bUjFXtrUyVjr0IG0D2DTC8pnAjQlhEg3IMPS5W/ptLxS/LbOlCDF4TGJyne
XgBZKTGZFQzdsuZtX43ZcHS1LFOKE2bgF6oVMV/h+B8OHNoeMrIulBwjPC5OVQp4EmnBwFB9fMZ1
/jdGyXMRYE3B6kUYYxIA5PhtMuFvZg3VJuOsXe1i0NXaWRDA8BqWgdymGD8JX2dn+gVSefYYHmeB
1NkEP7KtyjJb2OfbNQzE6XP4mTrFz5C1pbexfY35OxCJydHBBVbr2oaG+y6DcWGqp5N8uJQFy1Xr
l+ighsAhjbvD3OQ6cd04JZHlhKvBIynyknbOPQXBEmhVqaHHowV6YW8AF69evwSpjjiQG7n01znM
J0UWuTCSJIk+g5sMRqh1teyflZQnMvGsqcFGWd/hOqAl0SCv8FI39kU8TP/cwFzA4zHnpzhgMT3u
W0p7JE1oZp9MRthYG9WDbLjervj8Ob3FBrEBhVjv/NtG9vuZ/y8OVyCrTJUAiPVjzj+g6hR0ML03
CWT4QQhN2aScEv7aN0v0LuEUm9ex0u7j2FDHbSHYU46yXloB9ais6aF0NCS/C1vIPMUrdppB1PZt
OeeN/ups4EDUzlrEKB+DhlcHUcgZAH90AZmVqOrBERIItbMMcNE/DPMtWLu59tK8Gs1RwnY251VR
ycwbIr9l5VpqZVc/1/3nr+dR/ngh9kZP7Wr0yDhZXc9WflswFO6fe47UDKhkKLQiLWkBOoV4gZwv
vzyi9o8zaxnI6y9+xyFNZlclcjt0h9leMhXxUQaool/tGvK8DMQsXF1yemQHS/o/bu4mrVN/0GoW
cwsT6ovwOgyaOUKeBTT5F2TFZ1CJjtTfChalAtOWxxCIHjJili+tNdhqmLIF15riwl21JU7pbxaZ
XxY5fBfqALz/4Zi6q1QqTpFqkKbsjo/dPfbrMyE5gmUlyzcnfRy6rSUuNHZF1bzXG9zuybC+7yN9
/ue8CHGyGqc5OLpwDWvrqq0tirSDwGb0IOi69kfYsbreI9NULDR/JWscpgi5XTuO/72V5lgf2j7j
fbv8CjFn/QQmR3QHCoqO0DIygszwLpZEKIn0hU+2ihpiisX9+PpZ36O3LuIQCxYY7Faz5hb8ogga
TTjU2/cm15604JmkE7zj/b/WcqgG75H5gNBaB4R2pRrYKlbPZLz9xRJYFKGTThLXgbvAhufsY5iz
LVcfTT7/797djg7+oPxC1JkZwa92d50Jufiht4YQcSHDjKWJm+CKnjMJJSTCPjUKO34hcMseD7Mo
IpQmqWidiIpEuB8nv1LS0NTtOuW+q1JWM/N1HzniTdJ72Jwi+Z27xGa/vai9eCHLiHBmO1XBzjmr
WZpbY8CurRvftn2fJaeJ6wPakotRH37AUjwJNtj749r+6SAN74OmVQaPgemSictpEsURP40ySlDZ
RCH6a/1HZ/F25Y4yvsUBr+wcwskTPMVRJEUIBrPdHsjQlSUVE7tJULiK2hNocAOHnVqaaIkK1hKj
IlvTWIts/PfUAoEeMO/2suVxc9xLdhRSYNZBUNnANBnJIq1psVbg14B8kHgvojKwPNO54tgZd6mA
D9pk5+vQDZe9tmgSPzEVmpri195Zxb1/zADBte0unYZSyC2rD/mUAmjm5JnSSd3b5i8sU4RK79GH
E1s1hoIpPP0caBjddrPjVllZ9XDXF4DQdAxRMJwY56X5ACAHD7U47LUyvpwb5/nKwH7Dh9v4xS3H
OBSRIyoSFHEzd72uUefss9cW9eLp1dluW1ZrL1I5JF7v6Gq/NRmEDPTu/vdTdDsu6qUckIId8ZBC
A6KY/5iyfsBacuKoAP+pGPVlLXMiorJSPyL0U127WfNpLqzeDedD1fMPcGO80m7nmmQ65M9Vwdn7
HgutrD7t/l2jSHRL5RCDh2ALc/lHD4hNkqLEtngx42EUmGxhgAgWhDNJnsUEIot+1821CrkL+aSt
hFqIQHCPTZY0UG+LhLmCMCon3xy67a5rqu/kBrEsmRX+plZYZVQNKfAlDB0nEuOOr5KwKLKoZ6c/
hnL9JUp1y2bSQFQFhu0jgx+2VxV9xzrXsdriszGqm9Zfv9/8HqWlZ4i0LZu8ijRu7na5jNLZ2VKL
wiPuJNF8F1AgTDLCYIWbTNFUrkuhlGJt70upUsw7ZEqc3h/WJdbgd+pLRANjSA5mhnofnndcntae
6ajFfRbm1DbKoOCo8sDjytWKWSbVCV1oHdZcP6Vg9AhCetpk0VjttSvW0k4hzVLfFegYGsjyhWJG
XNJtl4K93Vp0sj5xfbPb5h9i2Ba5yswAlWgp6pg6ZryMj1GT7/iVbV4RKPVjXibYuO89oE/mOUvi
VOpPSNHJI0gNssj+EUzhU+yGwtlZ/rsWkY6Kl8mddHBB90G/58j3r3p/OspRjP72PDKi/njzO5VT
kpdPYrRvvn9GtLpQUgXJJKhYOg69YtGA6xyX4ODHawRp1voTpvQdgZJo/UT12t1BJck/c2X+FH64
MRiIcGCv1ZjMQci9NC5GglJfdUjaSgMEl0tCCD14Y5kFSLQl7q1IPYvGXMwUwzPS1t3XJe71LhW1
IUtbwutRUTi5OcZcUyR4o+8e+WrnSmMgV1Vnf6h6TPOZ/n72HyzJ0ddIFVYf3RYEZZ0XWVfJtDmy
0nhe6bkKzAJ1PzbMr+Vl0+A91N1ih9zQ2YR8Inf6LlZ+AZcpFEhjOY76CdIVaF0RgXXqcpmWu+Gj
rDOAwteYygzpIm5C+43vBwos4d4xrF8qe3i1CcUIUQtKv/Uls5O6788aUbCvk0rj5GBsRTg8iLez
uCOtiPvwYxq2w9iLppJsSV5l2TYZgqGEOLhORIXCTxsr0P7dkqd87nFw9NQp96amE/BBvNH0S/zk
uFrUdsrbhv6Ajg0kBbMmjfIybgO0vNepZTbZhGqQEWE12IcbiydGglwKY04Y9IB516SZm/Il7sRU
Wbr71iRNcgDfmcYeemHk7VIBo6k2jdSh6alvxyRq7yzuPzZk+H5OHi9gxIRxraTX0ojFNEjuXrPC
7c/tSEhnXu7hOao2t2jOni9WrPAfdDAK3naxvC6lDIk+d5QoAkEbhlgxN8OApGwLFOQNwlfuOCYr
NeHRp+/0/VJdoYzBT0/1CVlV1JAh4JsdMIirjGZooORGZrh3AkDBX5pqjNFV56/RSX2qaIH27w3A
aUe7p/0gO0f9+akjjYIHQJwrob089N3Z96I1mfIrCBAPzJ+MEpDpeA0+4FqUU11ry4tfS2Jd5zlJ
ulJ3OEpugx6omXsp6FCi84hOaHca0MJxocZMC8lsbxFgwcHKy4plizmndBbChXkjGBrt6YRPp7Zh
5a+l/hVh11gcEaepqZktLU4NdejXQpMtH8qbRVKj8x0OHqycusxfx6KBV5TJYXdWZaTlOKb3b1YM
8yYqKlr5DJ0pD43XWFUs5UeTF/B1e6I0e8c9CA7IMbaOzDj9n/7UHAlcVJ1DopaAxy2EYrxKR/Am
wg3RrbKOtR8Rk+DPtUTluvq3VCmXheh0LDe1QpmbOb6bc00oa8g00Krf/9BOlcAJgTmdWs8ciXr5
aahPv/2xhMdUla/IvilDyUiASltotTlAF30dDBOcNQDT6C/qkO4hI9sLEyg3++sQCvQuKnAA+LMb
Gb3/nCaDSB3wJD4nltoehqFBU64REYT4gxhu/Ufkf/0uxTSLl7DMh46JGJAkbGXDW1bECSbESNE8
ZSxwAl7gVXn9qmljLMaY4DmXFVqJgoKAVXGjQsVJ+60nNA10oKr7sFhhFJ9JY6c4e4ASG+tXF6JQ
F3NA2yM9ZRCdPwaasWMSPmm9iSdFcQjcri5ajgeAyk7dT067kaoDOabOFczutDYAxBLxfesvoZXc
Euf7c+vVKQQlBpFuLFR6CS+3N21cPtPn20mUa7EnJKfuhNsj0pwFEGVHzoz2n8XvmzRERysZlqUf
/FjZSOtbruiwVpn1D6kNpqA5hBhzlW6WlFmeSx65+61Jya/wlKwoItBafCoqoAZdIHc9704Z0kg6
IXZ5DNjM9rJmG1bnCiDFp7YcWLH+aWyYSlLs7rAbWX1gI1ICGAflNuf7vgxrpn55+5goVuwqBe3Y
pGEdtYi6Bl2IqfwvFqe4SzD0ERFzo4VypBUb4f4tw7akJpeub/SMyHzYZyGnPeFh8g2lxfZ/ugxA
nxLYBU35vwP7b5KRe0qLSahQVe7YKM+vXu9d2hUoighmoVkUqCcoV9p0TQFI/GIiG4tbu0djJDa4
J7D4qPgjyv21PeRi5fEFmC9IVgKx/GSRCWCue8s/oixXveiZsHCaPeHoC+GmUDq8fuje1be+6VuK
d37hQxD33U5U0WrFDeR0LekXeZdPoWPbK5BwEM5vvuH7qxgOFhxlT8irPunYK7xnpAKxAUvOAZLI
BuIwPaVYEIBsepNKBYejBOoFD/PhSSmDgHn7YB3u/dB3FRJDnvVNZjXCJgMCXT3T8lFFogqxPpKn
i5e9poKtX7IyjApTbQlwWqFQboJahfyhghyHUf3u6urvEb4y6jKLEId2MJGnpcGWK53t4m2EC2K7
wOD3yGc93DmddvQuML6ThMEUm4+gI/suI2L/RGuP+moLHitwrOknlqWEu83oNQisyQSgzdLqz9EQ
j8XtzU+4AS2F5yUaL0wgfvcRAViU19L8g/Dvfi9k/lAlF858KDKpA5zv5Cf9IxMiaVAdo6axtvNp
OLg9GV0jX8epADdnmtobjh1j1hkwWR6JN2PxQOIvJAiJHtJD/oq+lT/ssOLPhcKJA9UzdnpzTbS+
GMDjaE9qKjK0x6rYNfPYFjaXCfXSx1ponuQoY5nlw6E4ft3C7cXoykwhdDOdQTAD4b18L/tcs+zs
HiprjYkfABlHNOYWuMhLugpi/K7+TehezhUf4Lia809muxxqe8hzWfEtolJSDE9qJTGdayrqebr+
N3qYavtrRGkQcZ1jqVVSND2QD62sqMgY/inOuwhBmRFN1/fyMOvE7Msaci7VrU3+05/uZ6z8q3Xt
F/i/aUbIgXOzu0Px0YZq702Yj8b4hy16bbupeZjKtZnl4/OnfsT+V7yTS2+9AwAC8GjnB5NWaoiQ
hWckSngSQViG0v1xHlD3mIIE7F/9ugQ70qsvT/3tU2j+J1KlemGzrhj/LM4l3PtiWXN7BfJr/mLr
KDEG17eYWGyBmgJ5JCgxW2s2skJJmyZbdnLKYwRC1e1MkDnj08p7G85z7/+76pdOL8uOG1LnF6+/
SYHaUmHugRK3C6Y2Vi2mHg81krGycc1EH7Lbuu6R91IAOJolefOpWZadmuK48s2W8Aeadx+d+v5m
EXsl4kUuZkOgWTkdDeCYi0RMass0n5kyfMJmLU7gEGGo9WAB0Ls2CI5K6AVJbeIWBM6vJKtNQ4Ix
sslAR0DgikfxiN6GcdEvb/0m6lySUCm+at0yePGs/uWUVbCojBjadIcVhjspsIrwLorgyKSMDfg8
8odMn//Wvcy8lt8lhUZcaKufWQrXV2DGUhqyTS0YKNtvhjvJ0FrLABRWw78qQie+J32iYdSIERqS
tzlYeoRPLkI1ynXTWsd3oaeIMq8xvUtRdXckeiB3Z8HZTC2n625ND1iB5YqewzU5nKG2P70Z4aQ7
toSTuK0cdE4ZREo5v4p7+7y9/KalpmJ6NRxPbZrUHXpfzWNIir9YnXQOYYS99cpTIOw1fgLm8pZV
4ob8vkiSq8un3yVx9TyhXyiKb3FlD+In4qJpEysFF51yTj0WdGnAAoYDf54dLVTPPnqGU8dbKvnN
r2mSNCM1XjSrgVqdC5vfMei2nwIoWTHG1SVM30jJgU488kasEZlhECf2d2JDn26dRHwF/rWh+r2x
/VO5biuSa+5VqeXrOqzWPojXn3QcQxLetZ1uNYn9nspHXSTAc84YHoM7xoNsTQMXL0ngClqFrNEt
Ilxgjgj3JpsvRSJQ6rvtzOE5kqceHJl2RhnqV1Wk/e1w07bh7uFdm6PoQisMxJ76Tm2CFIRu/j1S
Ejnfm91GceEICAiS3PIghemNAb36Oulexrdon+IroZcMv8ICczYI2zc+T08VYW4QRbmcrfr4YAAJ
Xxm543yvUnSTqJq5NZ+TG4m1cmOj3iILQAn3XszCQbMGO1fVDud8f5KHpEzmx0Yzbxq18V2piIfw
ruGyIxIOrsNIwmQpp2AoOejrMp/bTOCevZOHk/m3hsEg3rHczekmUJmEoQIknc+VIaSV7nwXLczZ
rvUlwKFj+S7J9fAt9q0qvQWABHhyF+vy9GFXMdqbjgux/9qSxC7SivDLE1vOvKYMQj80I6NLpmBe
M7Tm2j69IGGF6cK/c7mUZyPo3R2CKXaY06MbAnutKbUZWCt5JMBnZjtyhKkMYk6wDxD4L2F5UBgG
Ty5cdVlN5k6LiI83JT+mYXOGJiB+EOMsgXk5UEfCc0eaU8F04ukIICh9ZJWfW7vcW53UPI8j5XEF
DzhaK7Cgi6H34j8RipfkMMyXqV9565kadnqOH2x998YevWoU1xYqlStuy8633C1WEM2asUaSkGmL
OalJi8S3DODVk7jg/DhQswZCNZhyYT2PHFEpP0MIXtPDhfseZWnul5rRXePl6kojIeLEjEConlJW
pwYsUNpx6E3CYtbgTVJJ6cwWjrxWp2SlxkZO1vprBF7o0XpUkj60CzVIJc6C8HOk78tRa5uWI6qw
XiYDEfC8V5DNFHH6mTQQ1kkBbg2uQKn3nsSIrLHBHLaeJ7ueHPlaJHbvsAsR4DxMxX+NZmZmw70R
GrmJ73N7xhfWo8KCYDnXkqmA1BpF/AciRV29UZFSt79HbeUN8EmS9RMdtRgm2RNxrVSlU6RaW9Mc
tTnERaUFd3cHMQAUFR/jDnGB+gIgdU0y/CXM1notxFB3zvM4R6fZEN0OYa6QRBjIm2xIZHALhPtZ
k0T1sjWEdNTAnTJSyBcgB2w7NQ94ao04h9zTp/AqFiz7D0dIQjKqV7eDvK/T9w2a02zBpuyh82lr
UpqmbhZFGcF7QuPv2qVE1NSGdZEDpbVgHgK5XF8aRIqC5/UiJj8l7cSpqbqb8UmaeVQ34A6HkEih
T5IdieNirZx+YPElRi8OnpfZ+yygZhcLXfzEa/9Ho0vGjgx1yzeCzdlSrsSAC0rHD8jakBGQI3ND
CgUHlcHRo1Uxj10i2Xq+IcchYzYBk6t6vM0wVLDcZ0l0i4YcCMe+/akMyOP1ytxGq7MKp1w9kFyi
mrUXJQAZSJtU3FBU4Xc2qIweZgl+mZbmmjQG5WQyzVJqtxNnb9sQssBKL9LNou2iNAzSc+iLoJc4
/e6HJJTVAPdn403Gc5vEp4W2hTdx1KzJ9sEks0/2zed2CLradMvOlb8FE5mzh2cyw2Ha4Lnk/qy+
DhD8PigrFxmWEwOuHE2CaLWVzP5B7Blt0+h3RVhDx5Zkvggv6ZtKgzfh1Xh81teaXVcsrlyj7FRn
zop2kji4/OtK27VFPHp9NxSXmDQCynd790UasBdAenz7v2e+BNrmBb5BrkLj7Mo0ppgj8nDxHA4v
6E4ncGTtp8RM9CzNFjva8pELwSU7hjQ/DY0tBPHCwqWzdQngFPT1hj05Na3/1y87roHzQ3dHVvAo
TbqhKheC6wghAFNQvk5+Y7QXhNrm+eRAAM/SbmDosQ2VeyF9exH6ub8MmBQ+G+Nm1TDS38tFtVZN
IcEBeTqjUB6zOg+42K41o/RtNYYRpOM2ZhU3Y5FbUixPYqYqn2UP+qckCT7ZD0KsH3ZyMFfgR8z3
Ryl8auXr1+gU/+eSQIpiAPMHyqeYDkmtuSvcTYF4SLyiBbTmmvA8DS2vXoV4CCafNVom/Y8DOMTE
mlWIk0s7nsaygfj2ubuMUzCKKE0lDuqXjEGtqSwK/uZF9M+rWOPv6m3PclgC53uxHRDBrj9bSGZq
uPhEH0EuU8rF9m+cAotS0peRbBtxrBOb3aFgvhOE3mvLITVOTYFTts1bsEZxBi25WuXxRcHgAFht
Nf8qaW2gVsBX43s9HuV3Ij4v+kurtHXM7MHdg1a2cUQ5xlL6ZBlq7+nkhOABnEVq4aNDTitD0HlI
P+XtJtc+1XpHgr/0V9jYEamL5R4Q6L4wrUeRpUACO3Ch3nJi95FdTExf+QSNAQsVZ9G00vJUTM+d
wZwFrkCrn0gaYqXJm6QCHuAXAzpRyVADa9mbM3ueD5Qx2lkhsVhCdpwMd/mpOgFQoyr+GvnO2UBN
hZhxPG6x+P8zaL+TTkyTzLe3LEZi/TtGWAoYlnD0EcEn6IPR1+ZaRpDwdRti6NhvyInKgH2KWL7Z
HchqjXIKI8lm+E1Q4uvVi17lhdAnE0M9ZAU+IvScBOJzB4113OZZxxohk+ljXspBg14T3jveH2UF
qiGFi9EQpa+ti760cemN+oz0EEHSD4KY8pOhJ6ZdssdB8sIz1ODrb8/zjQAfrwTqYTV3qRUlnHfM
+2B0IvWH2Tfio7gzCpZOjWvg+ElgwO7VFJpZrp0pWSU/E/3kDkuBhjfIpv5OWO9omJtWcrtG5ARs
XrrTu5PHogtEujPOEXDNdRjqTIt+6X44OZj9uhWwdVD6R/vuBcCu27dpOp/jouUMicMRWGla0Juf
rG4flJA4/sMCSD1A0D/W6hJc3n24KkbUSnIdlwCY5zpilolHLvSIerrMb4vl0rY18NbFlXVCAvCL
+Qcf5J64RgWfQZV7mUSneg4LP8WAiPjdhoBKj6Zh1vsJmKW409QYa/RggFweBVkyXn/qhuGwJ2RB
Y7e5rJD/bqiS6cMHvGotQzTIBVg3wnBo465LWUI3YaK07b6Ofr32lrQAPr5PLHLSSGF+S017AlXo
QWOFkJ1r4k5AQ3qden7bygN9cjtogYfv549LTK2wKGO2VCpEfHpa3BH8NtwedwSSgKdDlW2EFeRq
7fyRKH5EXWHR0wwM0JTWv0mwuw/91McXdJ1TB0xNoeMSzwUUNLnW7tO0X/fpcmM3tWWotX2aoD/f
w1LF1I6E1HmW8vfBiv1DksXsLwFUI2RQrSt55Bpb0mvVIPWj55JVCR17IR3IVdcSl3PHJkCIGwdM
6NHzYtVOuLtJjN3bxgDK17Bunvb4YHsmuomQ3w93yYNrD1vvEhEEHlB5lFRtYr1wr55InnOXOEzg
2e2l2rkKxSQf/aUjs9lgkplhq3jC32fgdixHfky/wwIaKBMXknSR05NlG94XR5O9gfKq1fcekkaw
yFxiZaUH7NchLp4CE6nWNe7IaKZgfSxtlZYHuj7dGWCv7Eq/x4mR4NjoK6TxLPYhs/Fl4PZ8ddXk
3wAuGoVuWDST/kIrcLoyz0X5PxYp8RtSJvsMzhaeod/ua0T9tlXaLFPZQetg6bSb6EjPQr8GbOwU
CLLNLX/GQMzVuovzbjweOTOxwI4o11CzFKRq51bX4IjBQKTdy3NqF7eXJlqE9KEPAzzUQQ2aZhWS
Pysid5X7b9J1YvXxdhZBU1pA88lVDidP5SVuqrhh5Wd0NJlIIUG5GMVVTrQzjdsI2MKxoyxhz0F0
ZV9/5hfG2RGBoRkukGsTHtYtXkFqn6kiazLoLw19yjf1l12mTLM4an/7s0G1Hlt5z2rsdumP9Tpl
AFkgNKVXTOfgm4Y2b466VPFrpe6nA0p7NE5CZ/lC1ptQ2of9apSg4IUXuwEMkMVRtQ5av3gvAP9q
Ng7l5Tc6nZ6xr6B74/r+MqZL3ufVX3QgDLoxFlRHOkz4cDDnk6qdEQHtjnnGGIRWT5uigWG3LnCx
dwQZl1T+nZcQmKkhOjDHIyVzJhQXm9UbMVSC0KlvtE1mwzbMPQFlG3oNe55HsoFZnvhDI05y4OQY
efIad/8oTjc8ppcZyjNIoCZUO1OZ4iWBNqC0vIQUdzYo0UGsShP7qnKPRiprsgAVFqMe34P9zV4V
rYQNGDkGt/L7mFp8IXsewcr7Csa/kg3hYJItu01zkIW7lGr5mHXG2Qs5PabMUaEiDMf8qi7hLyli
u1p91sDh2uQ48MxEo0E2QkDahGfjZIT4/MB6Ap8Hgb7kdvQwQDqKSatsDFJN4xnGodsZzsCLiaND
6y9O362Ii6qauGadw5hn/0n78dbGEaJaxGS2kjB2NsOt81j97T7GiGY7nRAxUoX1bCHZW1iw0wLr
DyoptLazNlBYg22uc14pEUp9BCJy3A5rtQtRu7jX+TdJumIcjJjb6islmqDUkX0BpFMX5M5Lm7oi
XF5gP4UuPD+Po5iW4qHjmmDhRdxbjZFqNWnAyzWeVrNLHzIie5wGdeupnRVNbVdJJdzXDktJcfc2
KrfITCNnhSak837CMRp5xfDN18mWSJIjTfPD/UnWZNyKC6B8pTIZqj3gqtj8kMss25suw1wVTnyq
6Npy6T4p3wDXFj65y2I9jtYvt2IaRxyXzZwIyYrzJrCNMYiaBRUhvckaxT87H/e2dpFryC8LjXp2
ZOoKVUiEsYsG2tHhvLoForc4iPOJlnSsA1OiNPqQPkUAPfw7TE9+LXVIGxw3uDWGkEYNafz0RjHi
Bqb28g5GW1XSCqc3QTu6nXAH59UgTTh07udv/GSZlPIbgLfOyjW4YBFzRiUSyUn8mnWqnEHQBlCd
jW8nLcmYNtlPIfEmGBddeKjBtHJMLskkNQcGdb0fOHuF7hCaQyZr+Z9lty5e556AKIRQfRXdagC/
m3NE+ZiW6njcBKgGoZarp6H0Xx8qqdlcHGFJk0bA3VCjnQp82RoajrTWhqLZJgmIasShbXmcW5Qf
Qry1DyyUAW/dXnatPKhcuJGeh/XGJgNLw+2xZ+Ay8T4lngUDnZTixdGCiYmEhf4zy1Z5gSi3Xk2D
79avLeSlKKqBfJcdtnaHm6e7BMIEPeB3VeSO6mrRa5x9rzBYQaj6qkBZ9Pc+3UsJiAN2rDaw3pIq
9W4XpTCJF94UEKxJLuKp7Hg6wyaNvejp2VEEzP9/iBG/0b2JAWgNU6iN+RnouX9r73sMCX8pGUPu
cbZ7EhIIIfcW6C9JhVup/3ZbQ4bzfeFPkClCQsO4gHIT/ENIhSaxhCMciMt8ZhWwZK4PpViiWANz
yks0nt80EkNrs8D26GRKKAB+YnJGP1NDw0HyQyAqOJyTIa95st5cpOnmlG0kEAcdDvH5oPmMs8ez
q1JmHwIBf9d7rDPyY0vHaqV409y9bP0fcipwgTfFiBrMBi2C1nAL0HMGjzLRiBFXnfe3DoaBndbe
KP/VGeskrXGJ05VmRCXf7Fbi1MOYmM+12OVc4H9wCoEqOak7ne6gi39c8mbJXzWM0/owO/X3O9qm
pAed5POeQRp3KD9ioZnQJrJSUgGKoonboJQZ+oMZ/Go2RwVc60CZJd3g4XM/6JEfAklR3CbheRuJ
fixlLnJzaUOeqenQoIHPshID+FLNCPsVjbWA3k5JFA9ts9Mlzp9NOyNQD6kDshwRZf0Ao53yncYM
Nq1AtDHS9T76TCwzGdP2311lUX4QeV9TKIXvfaAwH6hHZQprNCPXW5zUBaCghwNnNYXoJmRAghQJ
qiboOQKCqAayp3cmhyEEwqW4KIDYJWwgxa+dYbOuSNN2XbZJQeoSrQtIGl04nUQsHHZQX27f1XSU
s8EeGXgPaeIlfwVTRJzH5FKe/0QkrZFX7qmBUFmpN4UBZ9901K/bk0iF30AzmrHZfR5zdFYo71aD
Cmpfl8ZoJ8hQE+6KrO4qyMdSZ01kl3o+DBffdQ2tsfucSoy65AnffY71AF6v0dWaiNjUFZ/lzVYg
yriXuC6hloo619AgmiVDf1MNymAyXKDBPL6o8fFDePN4CgiiKGNjZAOm8CD4Lz5KGxyZ3Pm9JinC
bL0lBjLajfrMQXrixe8Uct1h2OdtB43JMYdIl1CehqNBP1F5ei5LplM2Ejx9ehPkLaQczYEYSXbN
ke2TN2SIXxIapJxhdaq+AMJp15818OKnkvwE3xeAX+1vA6nuGh85j4pqJ2qi1SdCe2U3Olmdc8+4
qwQ8XVrzHrx5/5tqWMgBR7SFZWebyA+8yB2uCoYg+r04JrJNbN5Kgcfw/VeLztd8WrZd5zDeckwV
cwODAnw6nPubJ1b0Qw/nK4lNNb95y90MHyAPe1ikwYQLGohgVKNdhyKY03jnVPNhcgoMqii3UFOx
z85vzVAzYUMUIjdJpT4174xfw+lyW+JWCFsGoex7GzxkLRqlLx9ZjBdx0+1ns8whzmC5Ou3Ytct+
uVNXNiSmK6AY7ZYlVqq5PiBJwrPf3Jep1YOsIQzGpgVWybEu96RXk1pPIvM1Cjm76Aln7VMyOXY8
yk+DDHlC4uDNQw/BkP/3oToD75yUM4TjofyAsxyewA16qkf1g0EF30+/gwXLlTBLsAVQsQWrkgn9
jI9JViklOmsKATYdNed+fW+kRP5zd3fCezROF740qGahPtbcu/+W+OUPK5XMj0hs8ViF8Vtv+Gi7
BOcS/Qe0yhS2qPd8aWVrhwtvscLY5Uyqks4zVGLAGTzIy6efFUce7VyfIVZYALt6nnTrdRsml4Cy
fuLyavlNjqHcvRtdw/F+WHgKVedhpD1waLRT0FIFxOzGuGKUWT0UfqTukkh4D3NKFDloasFQqte+
czvuUINpkBzJuwEpqc72xSIfPkEC3huNbS+rbuZlrAF1fQEVhZLR24sBpiYF88i+xlcyVHFW24eT
txrMbnYxY6sXSXEPsRmL8C3/dcW/aHwiumty65L3rUpSGnpMnKiumVUaVUZqFsjPy3T8uqUXHZSJ
Ui7Fg7VeXTP1MEE/mOj+vKcTOhFnCr4ok3xqrfvoeqfvZpNfFcTSjMbYK0WJHu2xkCPH4S/2UTlW
v0HRjzZIXoDap7VdVqvxC7wIDZ65t3lXdJR0YKAuyDYgHanU6zOPDGwKvqcSwiO9St6qEmM8SSgu
vNW/KTqoj+7shtPKiHu0AMzUKK25ZqvsCNIa52cNFJbdu/bwA0LQYUVyAeC83RyTUf4AMqf8kt/C
Vaps01bAGhneYrkIkB3YiZDX/Q0SLnfz8mGfL0N2WLsmbi4eBYeOmi3tyupYGKFVaz9Bx41JR9d2
YGeaJJG3Mw1jlB67DSkUo0qPfl+MBcFIppNw2tBJvBwoXwxHRApyzvmfZLDFwSdmMbGb82kpcW+J
vq2AQKEmdCGCYf+/5ECvWP1R3auKiwLiMs/TUD/qVH2ft3lr/a50CkuiOlgBruho09a27YsGmM6J
0ZUEU2dGjF22eQKDmI2SbDpwSxPSPiSygH7ZFLHYV9Fz6ZznIT341Bu5OdYGLjNsp0BiZiu9bqrP
LRbdgN0vAhacuBWZ1UY2/G5Bn98clQouql83gt8scCgAX/BnLtD4BPk0a9TGnpPv0iv5ENgxHTOQ
2kpkyJrOS71rF+W9VrzXKwwn1YS7xz0f99LGYlvbZmcv0cNkBPt7YxAuFR1fhcDbVtbZ99so4r4j
y7gWUfz2vGERm842Sa4g5MdFCp6BNrxJ0CKiNjA6dIy6xLIjDTDv5QnYvIpK6gbFtBbiFNFXskMA
QmxuOuBI6mDtcmN4Rl5rhhivgkqI8flKGDrK6vNbRivdjeMxJVP6Ep8+fJCdQrIfR1iW7a5SSIUG
1IiW0ss7eznH7vfimtW3l7CbUjvDfPa4sLjsvpx8b1PNC5wHsllspK69MspERYrfuSQzeyWeNQ52
xQgYpLddR+gF5UkbvbSJsXas8uwLZNu8OBW9ltJexXpD8li+WECeaJ9LUV9rSP0NcVpVOiGMZ5lS
FZkyKiVPSLSYshJGJkf/PN2Xp3z7IU1NGKQs950RF44jDV9lcYSxYmCKahY2Av8bJOuv38klPxD/
NuF5l5cakFutqxgGBsUBDSLkHfX4jIeprF2pn6LGhI5hqXsfYbZ3uOW4QqH1BkTAsXr+0Zm+I8Vc
JGdPF6t1wvkx5m24rqKJZw/8/808VQ17N6UfA2bsBfc/xIKSGpnDWam3Y1oBrzma2QjraynInXVS
+Ub0rYUcMH3juj2PZ2B9Xl+NyuNIzInn+hKri/eNmfrvrBAV8yTl9dS7soSIeiPp2WAFKvFiW2eB
KF/kQFjMAtmPpKG2tThd2iKoFO/ljesJ59NAUlNUzxzJ/nWhrHvviwKtUDnak8viqqQSVvYF+yYg
gBr5B2dmrRz3WwHI2Dq7dqzgt3Ko+ydH5IcvnNWBhr3SQYyqSzTOfVw9GR8Id0npC9SLMRFiBYss
LL+xhjH86HfsIKO3NnNT9eTcNHlkD4un+OTrDiPIaukgIMnnmtOWwJi5E6p8CNrhqVuPn1G2VxLZ
EoZ8Jyj2S02MR5YyxrT1ejNXbCr8SXlUBEYP8u6pj8O8UxG+9BhJVYD5q5Do5FkW0uI5w/wDPCr1
ccL9m16R+v4mWdnGsE0IJX6GFlZ62kBbuiAJ3eTuZS1z7hqkvrGseD18bKnqknfpDM5aJperMk59
bXrwC0HWKyTCo9V562AYYmC/y7IKNyvFiukYRjfdvRk0YU6yiygzOZEjqFkEkejoyWzaH2XYQ1CZ
fXcbhSSAQmCx7MQiyZZRmuVQ955sRXkDLeK18JHlLDdws5ur6kagREXm5wMHpo8M7+iwy4zq8pgq
9q3vZP0/A3ctuSUTw1I4uCR0x4OxpsluNJxdMArgCqg81V2exBCdn8CiQZgG17flSmgtY2E40Yii
b1LBFYgQi+MNafBuqJppzb0ZT2Uhefjq/DGZ4G1aPHEqBTliN5W/B96oDmQHy5Ad867lUA7Q6yl/
rTRxCl2/9sG7j7W4TfkGdzR1M6xAX8p0ayhyjt6IdspCXuw+sNeRpfZ9Ds79egoNahhhbwGQ4hlj
6rn1a4uChSclqkKBEJkPVscgcTWEOXwaeRB8EHRi2DoWP9QG1WvK6HhvFxwf/Vo+1LZwPwpDA+2h
fGpf7jJNp4CgpXHN4nvAAcOh+lr/Mb/EMeVZRKmrKIi4YGbK+SLnSIuT99tctkFr6PgdYn+b6ipP
VuNjVVkASb6SCctenp0zKxeADFxAxA1p/RxWqWdwn2rVrEnYOYo4dnInngxp7ZrQsr3L9bNTnYcq
lXaZ1ykUJl0oedY11dj6blEZFIaVTdil4Iygw9mwbS33TI0cjzgqirOfa2X/igKuRMmE2Cgihap1
eAABgXe07ELz0QJdWXwg52gN59qdhR+YHYjdGenuGIBa6HyZpV/NMOiisyZ3qYOu6eKh685x1CjH
nmLOTUQEr8ErBsJ/VnsrCB/ykuqGHhoOFb+/3JEOZM6W4rEGYqQAgez1HFLKNwPNko+fFnQNObT+
GBhlmkKZgiFt3zVgf2As3TbE4gi/hoIxUSkvACdMPxl73B3f4HYKwMtJwCDoPMtQ4LcL0NhS1b4M
3EmhWWXdlr/HgosR4oJJnPIRPOdYu+inKKhzyS1wXhWlFdMB0wRLZGJaLCkg8Ln1tO2Vz0sBos9g
E0AiXYKlm3Ox9k/+6K65z54uZO/TSQw1D4W0ZaZbl7p1g7dhcqUjFhSDK4MrYvA9CpFYxBuH/9Sg
mEP/Y0X0tXk7nO0PjwvtTHn8+LR2D5UHD+e0WmpI6yLJatc727YKYLXNY1OgOPxcIDLsdR6Vz4Z6
IyLnm+4L3Fr3fD4RoZ6Dy3e7fA6j1b/KSUnS72ddUp5nXSxZjNCWehDlajgZeR8ULVmOOS0YArpX
6LblfmAecyXuTIYenjoYeuPLglX2JSgsLQDnL98VpkdpyaQbZemBRBDgKQwCmP/R8+xhOLaavbYT
+LLJ2D/xQaKbVz+abXmsIKUSKUJwEl3cegeLFijt82Dx6LC9G5e+T/2m0aMKNtD84sSuzrK8I1tI
3SuxyZqGrJ7p9t5YU9bE8XiWQMfJDj/OrfvAnmZYHbroixSmWJNxTAhwzV2s5wCEsfwLn3XJYcC5
DqURKHd2GHo9nCTszpbQMMtwypFX5xGd17uH23vTQmqdQJOSwnXR1679dSIt3eNZepBJ95qteVkP
wCy334KOK8I4pyRhKjHvjryFTKoL3ZIDHfmDdJSAislyMFiJzmQXzgHjTScjzj9vsw4vCFMtzrs6
rm+nr+tOIOzL8L9hqdsMKjSYZyfpvk/EIsVCQkn/fdsGbmqYJ1/IHHg89f56r78HU4G92Se0G/7D
+atHctdrhiWso1joEhBpplQF509vMoePe23YoF1feeznl5MJepN6RbbYSblRV/eLHAGIYNXgDbbM
+wLsSdROu6briXCEIGXjuUwpKTq4lVhg22vYEKyitSRyM8xIFa5FU/zBSw+3eR6eDvfea1iVUOxa
yw8z5BInF4POFJzURvu9IIgDZkjZ6GFbX8oexCqO4WqkZ2NCEvFg68B2HO4tBJPZemFRaBwoFZ9G
HZicTZHsJnh0Lb/xwZjUd0diY/Iq3thWg+VHvpd0NNk8PlwuOr4Phq/i9ZB1n7TmbuJPxTfU6WOd
6KKSa9u2TFKYiWWwwbtrOsyMBsWrlaxTtqtV377jsjSwyknjjq3EdNwdm/dwDYMybCsQHJlNzWLw
U9ZED+WQe7w2e8hO8MZWxY1VJ6A4WfBjGRCEsbmU1S+6237Ihvjpq1Dj7u3Rlk7s4i+DKtDIntI/
pxvn8aE3cNz2rltU9m7u0ZxfE3E6jLoijsen/JHIxl8jBxy4wE/avHY5kswUUqgfAj1syr+cNy/H
M7I0DLiYNbDyRksYyAmZkIW/ifJxFLWaUb5bnxE9GNxBM77/PT448yziUdug4SQjBb7oKZwUUjXx
W9WJYxJNkC1XjN2zKyegjtihCNQK96651JxoTT4Fp/6uAv7PvBX7b+lk1NDij7X2x3RrP50aDHnM
AyLWAHpBCtlECwPJWQ2eU7oRB1ARTUmE9hhI30A+HHSd0oJBz5pvWHGBun/4TOAFmVUCA8WsmLna
bNPIQWb4covCui4mWH08HiYVzcbWxg7xxvPtFcsP9BRqReNtQ3DSCoLYiSqfPrUGDpo1iG0cWSiH
M6vRwNYtpSn4dyvj1tpKfoop3AyEMuykq+e4IGoHwMg3EyljQ4FNjYZKsR4w9cEP+T83HqQp2vD0
dP/ORFhJGXPyFLrNA/gxR5G/aRKLZYpemgQkBrmpcbZiARLL4Hx5bTm2svC0t3Mau5gwLadBXB3a
HtkIH4pQSaLmrKoj/jwdira7JM+oMb92tNZaiHGsAyTF3U7EWoBjbGr2AdfVq6/HlH73i5QGLBIz
NqDcVvaawD6+qrtP7RTXqPOyjHdkWHPCBxd3XzHj1/F+QJti200jVTJpJV+qNBRdcxrsXG12i79u
asIiUBxA7wdnS+nRT276B8MS6ySikTggI3hHFIOjApaSaiWn2sCjYyVQtn/6Wf3eX0AJxsFwl/O+
joWGHO53Z9VDI5Fq1dSmqKE93uYzfz8a4svVeD84Gh4C9rtxadUcA4CCWrkIoGSUfn9F33roBrb8
KihQW8Iga/5OqqBBNa7NCLjzCwRQOgHbhuXwnlBPwmT7zYYZVUfX50c/vApktJikfLDKNU2qZqsz
78aqDrh/dJsKnhMACadszuzkQ0kmqqghV/AuCLZpqV/dJ/J9da7N2+fKFXEY8HmxbiiTmyEaNrrb
lL9tn3BJpER3BdR7CtcnwuFXHerBDWFUW5Gt8P00QKuWDe9eh4csCFpX494kbGeMgjL4MPCT3nKH
mIxHD+olFHArZAD3wH1yH871TcvRY7Nd3/9kYkHYfNpEeeJpgpIkWJiLn2iO1wFQwh50vrhmFQEl
7MiXMEL6VguJTm4Nj4vFf+ymPpyTJbCy/xtMNxd9tKXODhRbCYq8kiZ3ZXqwOuh0NqxR4eMoB8cU
YW6/pV1Fo5CceL6SBBJdHQgYWTpn0cTOxBiyeDr5BhwydxShGlCVWufTy+rWzRAXmetk1+p6wUFD
6dIkMguxkqXvGGbzKi+9EeauMX4kXiYfIpd0mKOnsHJzwzn4KhY3jA3sOQlfpaLNvjvdIInKTGVo
Kt7ecA7M1/1Fq2R57bqUfNw66g5oiWi3SzU3Bs1YZ5y/+NUtK+V9dvLkWlUHXVNu5MOU2IePisVU
TkzZ/wcDrTHntlSq644RYG+dN/F7B75lazelEoimzp1tcQ98KL/jB1Vk45852ueuaOTkkLM8zMOR
GUK+hne8IpcSd5k4tq4qpXgBicLJCT8yqf6+sAm6/EHoBzKu9I11FPHHbd/tlSiLT6CCkPzKT4zb
d0BjC28bu2CSTMJ6QqpLUjm4jjlxX7L1YDgtskcZW1oufCubHDeqnSqClAF1mGRjeQRQZ+RRnbJn
FJ8Hh/4vsY6YixZlyNsxQEG531Q82C9NY6Z2OW3JU0kN5sEsgxQFYthqguWj1yuTBD0UAOADVYi+
w4iP+w2vrNicsBWQCyzjAKDJS3sIbSC0XfuW9e8a66hG7k74+oHR06J2Zhs3fSqv+J7roMln1J53
RFD3zlCRmRFYnkCSAVxPBzBoAslpiNvpwErlOfP8m453eEipRWVhdIN8uQ2jks6qgMS5YPIr60/w
SEZlffPf6bBKBpHZ0Hi4ZkbhGOkZzI5PvQ6PxCshh7fFt7ToqvCcvmMVzf9mAT1zxxEWu1qtcEcO
tVjDJ5z95yTwo4jI4idyl0GmfvWRG6tpTxsF/jJT6AIwvBH6nKBH2NbWMUCSjqUH8sKoYHz7yNL8
+BNtGaiK2aBrgHxLSzc9bJmkq8yUwIUewWl5YE8bKOVW6Y7sgs+sNDG74PgFyWLvc1a4rV6EG32p
3zaQed9m51qhTYVO/1I6aNTmGk+6pgBoKkHIFbGjjDq80aG6zztX2Y7TBX8+F6DhyyLKHU4AVUUD
t+6MMDwdmIgrKZeNmi+ZPHtV+VvgEq0y02xPZmCS0LeqUC08uMuuBmN+U+GsqrPWNyBSMIV5BGAX
voJ9lm7qqBNy3dsEz6pkVfz0aLOogcpNykgq3CLkvORhn6vtgwWq6MhGVuwzwAO61U3eCfvioQxf
55EXPKKZHMqrs5IYc76SjXf2+69Te5P19qV4H4adO7Of4A6rA4u7lJInHfuyDBw9K6OXvPSHXxau
S2VMK6jPOJWF7s6dSuvks4m5DkViY+dtK3t/26aI1XUeU07ijB1jc5FBekhPVdaeRHV/DoHePTuJ
dA84qC+pxBasT59IrMO9q+gvMDR6Bt443nWFWhXMouhgCOzVRjmx9HfcYVjuXdU7WrqLzKzJCYgj
e/Z0WAkMWV/qs7LRA4clS4xOK1fnsz8nNBD5wxQ+QsFyJhs8jwLekMS341Tjpt7kfFWqcbgngVyW
cYo07272GgPt2lqCYi2YK1zIlhvBIJvv+1ieNlZ0QwEZ00gy7qyHVR7GBJIqA7bGfeBo3RF9rx51
fmcFqs9vLQ7bJtFwU+sx56rdTLMmEQePLMAGdGRSaPcXgufE/uJjSHMKw1B60v8arxePZMJ+Sbe0
eLzLKqiBX2TAaCe3n5NgsxwnMNlEOCa4fRYc9cYwx2mlcYOwzb88oPYPYmKxW6pINjucV99+pQ+J
h97kIvEcOMK2esaAJuhFG+lAOBTmbOAkYvQSIWm3U56iSGbCvMQXssiTE/PYG8Zokw+lS6XxD3Hq
ehA/gE1oQOR0LagxOe4IjDn60eGfDHsBkSKQjavC/cS90AMv+1aCCAnn6cbEsZCYXDd1aCt70rUa
L99KY/WnkJhHmejbPgfA5csUtBylejlOIKlj3OZfJEiSQkt746KT6hhlYreBlzjKu9E//1RnQW1a
GvN9mj1G0H1d8wzNySWwS44CD+PhxMHPPcvjbrTGCtX0g0TqnYOl4scBhNeptqCpMQYx+qNhDUoB
wEF1JPyA+330ApheCP1y19M2xeuw2fcuSzM9oFnhyW77+jYTIOc1CViwtvg9u9479fXjnMpjkLFz
EvHA/KkMlKQ+j+OtNWyXwNmoeKK3dH+YphzooijT9LvNg3RtZLYcQAeboJUAw1TZMxBtfOYVpyS/
cXLEat3BocqklcTf4o43VB+5GpzlrfztSvV2U0f8CX+F83UlEJ3J7BQG7z125t3LZCdO91N8b+gv
+81pmB7dsNGvRmPH75mkc7+DHVKl2ZsGB5f/GALgqxGqUdV8SHxm/aLwxHPlvZXSABdoOg8UuIXu
DqLOc/HpD9UGd2hgA4tPi/RlOVOFXfu+C3fqXefsKJ8/7a3tybtmiedZ9dT5nA/Htqpu5EsK+LBl
vKCKMat6QO7HqOB2KQzy4/2IWMDke0G6kiTlqShjvtV9NUDszK+FaqUNVFhgSvRwG9jIB6+xkRH1
3/m2R7erm5JUJ+EjhN7//r7YKhcVHNEfrjETFByr8IapOpKlrzXgcUCEMTom+EkSNjnSKmhDOPRh
DRI+uQdsypRl5hP6xWN0rw/s5H2Wf3fK05d29wqvTXUl4JO8+AiSb8YaCVNMEpY9u5AnZZoa8Gwl
/S8kyDYtUQrkLDF7zgsl2Y8SbuKCoVyRWtHRiWrttrtM4oShu3igz1QNYg2nspgy8Ny+rnjeVOX8
Oq+teNiNITbwkg2oTvEFYjwwoU+GwDA7aj2Y8wQlZrA1sBPfwf64W+arbvTomzdHLmMU3m5pWm8j
hwvMNY0CjgVHiy/Ok16tCk4c8PovmgB/d1Z5GgcT+YBqkcobXT/789MLZFgO37/S7kfqs21J/P4e
BtnbJMHQhvaJmWYm1OWWsyiNlp4tL+LQzERZbiriu2sYX6/m8lpkiSDpQPYzFMB8PmXbxdhuDY9Y
5Bfq9gWKDPFMvrcwHWAV5unmbfqZzmqWJ4r3qI9jrLQsbr5bX9P/OoABHhTuqxobyyIG8/HRei6F
+OTMUIz26PFHaF4HFTVCKg7lq8XCdURJ15bZxWR74gM9yjvq3l79odN0GUVid3NqduFSHdOrFZzY
XpcIf/Ra42IZ65aJ0vMrnUyWhh6BrcB0YBiTLBdwKX+zru/++PZkbW84rrvqnYu0rawbKd/J86ju
OL8kNeE72PwttobUiHuiK2aMW+wgRP61w4UM2ychr6AOZW3osQ3Mu24P+v4YKNWzY1QQndwQwbXB
1iAzEsGK5cAF7SGGwk96em3+z9yzm8cOOE+yc3dcP2vlEUhRb07aIltMFZwlEIFof7LJdBZZpeCk
ZtyxdH1hmon2Q04U0grfs2keiqFYE5bp3Qid0to8t+0fO/PKbUAZNwq4Dtu3WOWeI4foEcDe6PLE
rpEzB+5zbifcBdhv6MmxQPjDjY2Z1d1IPcs9q8657MWhnfqELxsdSQZbNG/MFLpdf/KoismMkRKF
1nIg79AfACcpP5zhw9XA7ORXS4BpHKl4QKuvu1NwI4veP4HmwZZLfltGkZzoeW9NDyU5d1Qt6UF4
0lZ10XB5vwvfC4EQM0GsdE0Uy/zG6XLND0grAuxE18LxRSEXZHwWBAQOYM5t8Q3ZzjSUeBhwNxwt
wL0ss/yJDc2zeihsp10XzKpwf7FbOnGAzDv8pLLfoI3E+ijdSZ6cfqQQQyzVeUn3mmr2b3940kgt
X1AfEmLy+bm6Nj9byAbrU+a8VThQltUpfl7ebMfb3/34ZLJdt7UmU7znczxANSnNH+4BJI0WVZyE
Hkws+Vdavb/2itjJIBnReq1SjnQj7alERuEDetoI0/iHbZfv6Zjfhu3fr8YrWQ/x28cgL0W2JddB
YWjV0JkWmoy/82C71NPSjkloJPYYOjzSarm58dGNbaEJg6uw+9HEunxzg8fMwuFsLF0WSqnAEMUw
yKurIoeFEZROmyK6BYvS/qCM3/aCagAJcgv/Z3jcUAfxlxhesYiCwswPtBOa96xcSgcu5EF83QTl
XScRQtzMCM9ddEXaZMDOIXnY7iujw9uJ1gA4oDL9HIlDnZ7rF5w9G0d4bZNWuUieco0nCGSAOt2V
N+7J2BFjzNKPsqu1x34whow2mmdwGxLOYknMXaOrgz+iLKWpfC8Wrtr1a8ADCpGNj5JFltxX06LG
s+RvDnTG3RVHadPJFcBWFTYc0SsfbmKM4LHswy/Tx3yhxkGzPbUGejKVuIbEfePAHbY6xZGIXWOy
TOOPnC509N1+XxurKLT/U9LlFVQrMHjpljC02KXtk9NR+PiOeVg8UsK8+kP7TjUq9PAwIcrZIuAd
HYEf36bpojs7CnbRDHYVsPnSFqbW6SjODvfgjsVq0rUE4yne+Hjzzau+WYQbGx+AU+7xf3eSYQ9A
84gT474xzkdFRO8mFXDuloBqunzGvFmh/fgFfUBFWDkjE36fMG4KN2EH4z1htAHmlNDosAP0hhZF
a2JLQZ2J6xUlsFS93wv/bSFB4gL1i3RSkrAQHiFzFbRbWNzbw/ZpfaQCGNdTt5iSmRgmHQq+r1+h
AgeLMa6ttWFdMQTw7js5QxRZYOXDz7bnjlDAa8hYp747kac8T4niyWRDD/x9S3SC9FdZKxJZFVyu
tbfuICSUnUQDwLapzREBiOaRvRdPZqBKxSdkV47k7lUdDOpEFsLT9NTz4BdDng2yIvclh/Owrj7m
HPHWvTGfuHJisxkhszahfQhw32pPz7hD/Iju3CzCZPK+WyqdOct3mF1tVN8LrAMjMRm8JGAOWc3L
EPKf3BRSobEPUj7IgkbKaEMu5XAz7zDR+doqCApILorRcOm2X0PqixSIn41btJugF/jC/CvoS8cC
Lvo18hXShOn7HkixIAHgp5rlVcHcGVtVQiS6UBrbpgF46Ou8NJlGxvFgvrMSsp7hOxMha/7GN2yr
PpByV4uwuL+WglRk5KWBfhfCl8EoX+v9Rl4INj30sqUaMNfKYG9ryCGwwnPSQhacvL54KXwJXdJg
bGFC8t0h1HWRtbEbf6j4XNYoW3pCeJRjg0pDVZ1EVeVMEbFHWRgjynCy0zfP/oWFhD6J0toip/p5
CUfNFokJEzHO6G6fDf+UM4nz4v8IxeU0/OcTxUwSo/reSEnGmJJKACPAkB5bpZpMcPpcYM2zYAnl
ZBNeM33o5F+1uPyZpzEZpkjsh+v/L6hictz9nD1hekY4iKjC1JJ9GW9nKqtwUX+GF9EvxvN2Syxm
VJXYhLO7duh+6XdTrQssFVfmMOoTCSHlYtDYPeuELx9n4Wmrf8o7+8Ua4CmT5pQe0u+43MTo4PgT
dOojtshEdb99UctEfMStlFfxcwMBzXyA+2gZvLvKAbbRPLjMaeMWvnS5crc8AwopVmjWt85BhBD2
cggKdRob3Yy1WpebGk2sYWbOu9ApHql7lGWVeE0mF8Yc+PhtXNG7o01ctw2tJ4ax6gtPf6BafCrK
RUPJ/bZ3sadDnJH2aSGMofFYpRhXvH5hyJkm7Y0GmveevEy+/tO8iRvLA0GAbeGs1M3svnNC7YyD
kOW3Vfy2j0bFJrOjojpPGP6g/uLxcje8d2xUijMfrowF/FQaknhGImQT4EhWxcsS7Mp5D6efFV/8
LLJoIMWiPW0iYanWmkuCT5WSWmgheR9P/yq7oX/cxK/sGTFjjmyrX5ZbiMOdXSeHqO/cZWvVHpMh
BgrfAsbWFSMcEDu/kSuj7WDhmDg/RlpNom4j2r2CagkzHTUKhEwcscl8RmLdWHI4jaBHxj8Ugjmb
FHQ45bVca4qhWhYwOU56X5XeNMkXhAdHfhoIjzoTldFbQhZ2JNGn2fadCVu1OffguZF+PSD1wDY0
BXRz/8B0br1yiuTb/b2e7YcYeDruH/tDwuUVaqVeNI/p0uldSSmtYHnT2IPC2u8UM/y/4xo8tBcQ
85v6E1PGNelG5rpyTMHfr7iwERnwP+JgHm62Za6+uEUkHtpFjdFWBRQ/S/LVOhGiHYrCh4BY3fxA
CDJv/CIC42ZpzE56CvvPEXI0YN5dlLuBAnNwmWSENB/Rx67DSoovDSHiJzU3zY3BcAAxaUc18j+0
ZL273HhTWSEGb0mDxU7+JH6mxfEpc9sZlfud7pIyV4wy3CIpQVdrtdavAbZ0p9QLyKT4EBF+ppus
8g7KSvsIL3XKBu2nY+pYPPWjR8F5sf3vPnU/hcSr21IBV0Vh/FyFJb7G1qgoIJ4SNeBLQem3bO5P
NVanMvy1MvAN2+ZhfhhUg8A6EfvXn3LO8VPh9zZIdsPnRzB5onL94rJfxVRfgDvPbxY1vVHQ9ZY0
kavmmZuQ5iTXcSYHMcVorylDh1vQwy0udzT/MoLop1BQwEfO/Jy9GFR8XmxtfucUbdfKM/MjC973
l1453Z+Az0qcsEjHqxzfaQyyC6ysbt9t25ZnfICLvwYS5SiN6jMUsDMm7tjfagGmXJ8SRuKTcArJ
66Z4CdY5fdhtW7toAfEa5zybOrs1phGtP4tDx35Vgp4P3mzZTFfdFHComZUz8TIttvsb4hVp+zxp
7l2F15jvfY/HpASbUnPRSuut3YIeesVItkiJ2X6LarHfqyDYXJY2FDNWJKxj7sf6Foek+iHfjNZd
TYN3p0EmV7jlZJoQiNDeydY/Dt/dMp5XsTpMtTAoDsdR6N22WGCXQNUt2vFCW0D/lzVt0Ji11wx5
bS1tMV0EEB+j0vAChB2tPOmXgDUlYI1frghIYLI5fE5fWVlTe7tO9uUIN0AqGLKyUGIn63K816c4
FefEHCrrkbLBxx1XS627b2XuG8QLkD8kiwAWeYmIlKsu2COoXUY65BwvyHFwYV1q+/WUTOzWH+bj
lA6eTyzNnsZ7unzKo1/c4EEkFL8R7dDnVo9BzAXTFALzSXMNDtWh8KpkE/PFK1etKZ+vyl9BoWo4
/tjw5sV9exXkA4Bh/YPbigjrcyst5idUmUgtc0vA97p24wzOE31xa7z6d9R+Oja/5N2DVTrSB9W0
lkSYpKKfoLPsCUt7w+fkT/fNQUPd5tILIVW1l/CWIRWg3xhFjqySVvcgEmjzpyQ4iRt0KzI/WDvB
5rn4Vy3vR0kEqxr6W3zCBRnlDmRis5JGC5pGW8cTYxyPz69noqDhdGPWKcs2yi5xMnyoLvvXUymh
GptftmBDUMzUVPvehBs8vBn3nAAbNgw0VMMBCqRfTIpSqpHeluQgZuIcaSp3H+p5xMeLHpCPH0ju
wR+bYmLeQHoZJ1OMYyDr0mVWIRbNQORH1o210R5CeAFGpoKzs0uBv5Weyu96JqeTSKPsKjjKsMxx
BRI+FwQoxTpg8op46OATqzk7nzHKYZWvt3VyxrXLQ73Y6TVeA+nqATVaq2MSTKQgJ1XvKZETWE+x
ggjzhm6Pc7pvyfh/Ml0PMqvvPmZCnxibxYOmNh8AGE46YIBzX/DcxjQ2pZ3X9YZWns5YmHne5njP
w6xHOwvOi8o7o7vKq6ooXsDdRU0NqOsuPt85sesogPmt7GR1hC8BbR6Z4QowZlFS0UEs0QvPnpID
VsbK4xglYDVlLPfPHxkkZvYdN7rYo8U/y/eMjxw+cYg1lW2D/uUuK2EfuofCwMgwGrxfxL5fF8fI
Zf1b3aQD66nQxZ/VW0vOGuzwHjYMQWGaCLHg8uhHb+256sRfWxlfL3rmLL4oJxTkwCKGwD1GP9yc
2RAPt2SFBaCKDmM3zEepvjb8lMh3T5bDJBGSCluzbDJXwj0TiNtNpotJzGi9zl/QpI/rWQo2mIeC
AQihYcBOSrdQCRCHdBDv0tZoOOpJncV+WsgguqWraq/QvWP2rXDX2u7ujpeOaD4PaWch2YrMm/PZ
bF9/OmViE6P1SA9H4pzxMYlaaya36Tp/sl/Jwvr0iMCVMA3hEJX2V46lsOj9w85Ape0MiRgx96T+
Y1WkjzMB0GixIv9nMNPqJg3Ge5MRBJ7Qe+TL95+MyUrCpUboluEhHZ14y/M4n0d5xOE1Dta5eYH/
/SnYkdpDCqi9RmZ7Sv1lqgxrrLBzujrnkpWK1OJIsbatd2KHRDLyl/nym5bTYLVnzhDxPGlq3CUL
sn/5IwZU4+5xHhB4Z8aMtpBLCqMsZ3KIr6SjaDBm8SDQQ5Q5G5A7FO+ni+ST66jW3IdZJgD7D+Ok
T+xYGsuiB/x4mSoDXX7fVrTwkkuH39MYwelCcqutJ+R6WS0vNvKANajgbl3bKoh3/ghyq5KeUe51
HvvTPGdw2zw7NMSc2LEAKjQQ4qrBPqmc22fJl7kf4cnKTGXf+9txbn1j277KqbNhFEc72bbJK5zN
A3UUj+ipo/Uojv/NOUWS+eXUeh19BpF+UiPt8ZYddyGGfh/2Dm96sbBTujH0LVOYe8GvYQV8HuN0
LDERtf8jTvqWOjhQK7iNoGcTuVFoTsJ4S0/mlNSUdJwRsDGbCLYl0ic3uTGgvLOUWydmOdT/H2Vl
agU5Yj1je39R6kRZiGePEyTfbqFFjhE3xsH1hcTtNOE8rhALs/eefxulEFx4Y3aceH2NrWrtenEe
2d+ElO8J8TL+6iNiRYVRev/7skHcLmkgwEu58eZ7kwC6/pUyIVooEd8EoYNcoSEETApxTM16YHhh
YHVgCaX3MAN430/Qed/KTB1Ug1cx1IiwnxAPW8nI4V+Rv4hki8AHgWgjLd9ecsE4MeoxEPGI48Be
Ds01ocy4TA6szCe32TueZ1bVmXkRju7BsVoRk3vgSZGu+rI3OUIlkkmik9a+H4lH+EPP+2rOjtjJ
MEI0avgg7uilcG1bk10AmQOWYyy+FkNmMx5d2RITsWcuXDtQjaJLVc4cKaKEztcnFw/HEeJUlnuL
6r/G8NILQehuQmDnxj+ADVY0AT1J+4rQ+NUNhwmk2tVIcFjamTe5bch53636TNBB/FbFXzacp87T
Oh1/TCbNtYPj55Y4k+89EXwVylrsEc1zQxyu5ZoXrYBuM6I4mQLF8loyeFZSt/mJth0qkLitPD7F
oSmTZV7+mjG+oVKBceAVrPd5g4chpMIo3jlCxm7XQ5OAYptWuSSbibVHBISdFAHOpCnAcl79RviV
GWybf9Y7JRg0CH3BwlBEKEY04az1OL/uB/31LuRboAM3DGhDfrEpOhfHjM79qNw8vY4oBGLZhF8a
DhLTkyJFzBo3tRPv/UuTTn48BRz2TJyAfI8+fkWxymevBlyLAnuDEVfoR+CKOIEm0kn4eKju10Yo
8xjs4hs7+z500+/XLeBPWJYoymkW76OZjc0gc6DVaorYMVkWYewqU8zLoZur4eA1VOgVI2vWbm2y
KxoOQjdS52s/ssOy3rEEs3DgKUw3L9D/06eoVu5ovVR39iAAQOVMufF+YW8Z0pRTPrcngTMe+D2C
15SRMnr+47CuLP7bAWDBzK/rrDZjBiWZ6pp/tVMCQhtj1ukZA9bw3zYXHT4bc+kFSsWAF8Zb1eIr
ZQ9wzWeMfhpd9HWk7LX+D2EA7pcTdFEM0UO0OQUcfoLJhUX/MnDgHnZtoW58L9JgsGpPWxuPoOPU
nVEEWUkK/FjXhAEdT7PfNYXhG6u4oiEusamDtedjMGf/uuIKrwoN0E8S6iNj21hoV7Bn9PJWHR06
sltvW17Wni//3/7TGlDGtmz2v0MN6pFyVMoi7SMdONKaqKhLmXY1psdDYJb/dPiH0lwCegPepOfZ
FkKTasfo9AvJEgFWI0wrFojfgx1wxg+w1UGxs2FDxARq9mNIawnOEZIGx80OI7U4M2tTLv0/D2Fx
8i70O2DQQCDHHrOAems3s4sUYzr/xba3y9nOQK62uNH3TMKufvojnfyytrQZ6fB53LgFI09KWzpk
hZlGGUZWm3NLOeGYy51lfIeAxzNkRqKJQJ14I9iAb1cdVcQGwR7ZZaKNDLC1vwJ+hfDQYv4lQMCb
TXVhLf+xzN1rf+uUi2nn9cYqvx6rhou5+wDwRgIelcJGqlAsgTnp5t6YSTZInZO+lKFc3UFOw82j
Hk4pB58Jl+Rwf3AYr8Xj0uknQDW5lL1B+CA/TanmPNt+hr2VWcVIIGB+pJigI7uwhfelMsqoCIQL
5+vtwpxfhO4I9cUqQdiX0wGPo844yjwv6etg6q9MxMP8z42LXz9RtJ/50J6DklK/rlttuLCLFMtH
mJ0Zw/8Wlq/TOg63+pZCPWEDx3HVp3NOGIf7jtS9z1oX1180/udzWG1md75mGhWf/XaBK8MkB2wg
rv27+Rhm17DdgVtbM/nKB+AYLzBeaWe4uAmz0xOldPI/d+Uye7CpCnYp15ylA6wR6Aq6CvquSmi3
S4m6BbErAxM8ZKCRgrSX1tLQwqBkdSdDaGjM7myUVdD5Sbkui0plYgkdnTP+T2RPDfKkWQlK7AiF
kcvpdPmr1+Oc6fyTD2nWFQI+Kovd9sHH2ObeNpBg8CcahqPFqmMkOWuM2HdAWRC50mm6Q7kwjs1i
qDQujbw7LLIoVSbgyujW6HM9igIsvhBraRRmdzqwqGZpVABo/DWih+ERFBjg7kWgrDOuU6HD3eJn
8moIfCyBjWOQR4ejIOgFaVsQ/G3xYZeAHfvYHKw2543fZYvfrOHCGk4IBOl0EKl87HPuU5or7izE
ur0R5VHgHVoZDw2QOMpB91qYJihqXikGbMDwgqvAN7rP5YrVvQORxLECLx5c6bgF+bhZe6wzOM7h
ZTRaR5FZrD2psVBZpsknjOZfwKPU+PtAvYe9zZDkZq7iA7nm39R0uQWii2rfLCRkEZ6fkJEuREWb
ujPlomVtJ9ncsT/5+D2DzmWGBnUUcIuSbyeDFHsHwhySSMqL/Mpfxz7Rg7jcyMpFMbSfrJumXw3n
RNONBMYrq4jHRbRhHQDNJ7t9+/KNZ2Siwum/pDTgt6g9DgpyzzxJwwqFRU9BgRtlpsnQUJxkXYLH
OKhJ+7gMOSWh/jcD3oVnA3WkNx+HKVyFgMLipvtRPVR59t5c6d5Wu2X4SIPy7/ZlRcRzMTE49WH8
DvHoRg/RupKz1H4O3CHA4fH2d/zii3fPAuRD2yjf9fzXNmhk1qM1po5XuAj+5J9HeKRvISWv4BWM
5+ncIiHCayKK4RxJ4eObcdlpOU+JDCkHeN6y3lvH6/DO5nRMqGjIDNxO5YOmHBx8I64qB1/4cVOi
Fltyegt4o2OWelRKkXy/FBTPj/YCzZqG+s2rIMKvziBoxI3EilsJo8ycYVIzw0qi1i1FASAjZrvz
6VOsUhFL0DZSDN2+wTv0hdOicxNooonGC5VONH5GoRusejxbd/rJhbSpH1N703huJ0Njz0TAXrmJ
M1dRI9bdubtaXxfQdXCo0Y5ORZnWpPspV279fxn9nmAbIRpCq9DYYJgDwYVVIzXvQl4p9RMdSkGO
9yVlgYk0uPMAhg/d9Ue1l7V38q+UDj6xbZiGU3kDtWR/aybNznwdGMM+EAGkZxpol98IYHqVPtp6
Q1NkknUENDVDG3quIQziGBZOZqtywVYSIiE1ofPuSf3NfscAqEydCDvHLdtLZuLd2DakW2ZLGNuV
LLG6Hs3xJJzgN1qq+mSzxuC9h/nZFgmFY75QZ/9phViHU7ravWDJiIaY/YUlYxXs9zavGl7lrN5r
JDV6CSCG4H1i815XHm1vwPmXt82jx4pIQzJVlIUPrnJlHoJ/e8KzckDXyf2fsj2iBQWKPumIOfNt
4lL7yMAZyhswG33YL/MqfAJA4E3p2BqcBsSFaLfQOVfqcacg9v8zbhgsGU34zxLxxF1XprvOw34E
O4wkVwJPjeHRreYGQGquG+9uybocrvHwozgIeQvPF1btG8dCby/gdmaMKeAF4zoYEg5QgPeSB3FB
Squkc0vSOg9pESlBQRiUXqSLF7uIaoqqBncEH9b9uUOUwBMtnA6gOc5fX7w+ODa26749iIhTY2eK
RMExybOUgiUQVIs7RRxiJAfOc1R4XYCMfwvq2tt3yWN6HANLvqolZ8FWH5QDmzFo5aYZvwHUVIVh
LntOWxDzMZ/BLBzWxDE9oU6oIjZRMO9CVVwVHXeiusCjPq+vDUjsJZeVo0DDWraEIicyy1qT00LM
mG4M6sTzZ4R0XkcblN/KiniRUv3XZ+g0WNbg/PFy2sY62X0Ys9zthNCipJlGmY69hipJByaJKWJo
4KCglZBSeRuHXDHSwQ5Pf+tHRV6g41Hy7D1YKq4y6SO9K4IbE8qlSIKLAUO6Lt4kxDabqNFi4ELK
yWEZInUejfMGaUrpxqHKz5x+xVlUaNZ5aCTwD7q8NYZCsEKhJiUI2gHGYCaR1wQvCbYmsBZ/eZ/W
xoSHDqkiEqk53gVbgyZ6DcODFM1NbV+WYJBArhdG7WQMD4AAI91hkH+iJ6d/HJdq3RAG2KSxAroH
fJpseL1qZ0AqsVR4nmaBiLRLpCtD6gOEtj178Gm5+F4c01tPwh9eNyigGVcnO6ZOldLKY/uXvFH3
tb5lj/gT+YxinSsS7ppSwl1JKeZe4+r7DXBijrmPt/MdexGBTQTc7tbd269Do6ZBOuP8X95Q+K4M
Jj+KZtGZWn2xyMnVCVuf8v1Z4Gv2j6SPTVSb1qB5Pz+T1OGAso9LeRYY8Mum5M/DrDoIpnMAlmS7
Hfespw3y3rs3nAYzjkTkH60EydKr1RVMv89S5zn6BWjR8o1zhjTsmy9i4/1B0+56YwyRA1M3w45W
DFmesK/0CqA8DafA2HtZsSVn9FWWV5Ubh5PMMyWudIwWz6kevp+nGOcDhHCp8HBxluG9YWSEJHlz
z5RVbiDm5890I/uixq/fOIofceeNuQYxyoQ0YdOiRgvqzTqjVaFEZu5OiQuwl/vcfFX7zChjY4gU
9SZWbARa90JRbNEWDdjmpAnl8sHSooR82DzO5DaBfdrJs8I+cs32XnDefhoM4spMEzMkGowPDCk5
vvKjrmo80FjtibNRfPwC9wALxe2DYq/C4X52SU9CmthnO3i469q52wSmWdVpmR6xZR4v+CLLU81X
Ock2cZiqAzLOnE8L9WXxP2KmY/TL4Xh+oIFc7K0ZmOO9X4BHODwDMUctqbnjWxR5Hx5y4D6ad2xa
MZKXgswP7In8e6pNOmRX1DEr6PD7VUR1yd2p+r2w2siCqDzk0BH6WY1ht2aDz44hdxiCthx3ZuBh
mxVtR2GqR7bUhfD/lq8bxUU7yGgDL810NwdLPHFz6YC4l5sgB1YPtz08G9kzvwqMKsQnqEcMahx4
c9+xdAkB9yds9956AR7Ymi+dzIgCeI950r9na8sndEtppVfSMnI2x0LXb8NBkBiPTxRiDzMIAJLC
Bsj/McNOJhGJ4DDOz3hXPnlgXcpnhGMnyLBrkG01/IoCwyedDjpH97XApsUkZ1EA0TrWtfUdkZAi
m+hCIlilGmSAvlwGogCDlicGxgSN66ITVv0JMrpv1lIRM6bgofGqGFUfSzvXXYu6ka36hoYL2nSB
7ctY6IOI3eLupoH9a/3Z42jgLUkzswSik0sYM6FDTgQEiPmv6LNtuhbLDqzP3rW6k2mbRWvA8OmU
imarGYxIffGc19HAfzLhAshLsriDWVpiV6C9T52I10iw1bW2uwBFtQWLwGwZATce4mKaGYdQEDAn
lB/quVgiDuEwp+SXUz3odxiNWIGycEiAw3qieyEh2x9+0vAbkeqvhSyQZr9Tfjcqo8I1vcAY3Whr
ExJmmR9iI5Eg/2Yry15mKNI+n16LCW6oYwnfgMlZFkYlfVuxQqzV6HpbiceyMyePMAImW3gIIMJ4
5v/Drqs2uG8wL35frB7SXtAMY4JvjzQLYtjieU+dl/DOUWqIdM81RChnz0bZGqM4+MgmiS8v4ce4
22TtfetHewq4HIcLXI3/pTDJ3uTwVm1jMs6RFfbf9FJDm+lrSuucU4sWuQgkbjfaEYBMFGaAzMyZ
d9Pz3ieHL+v8W8W4quouqmlUUR4SCnAIsSweLSlMDS+SiSfTEFtl24A8BpNGSO2UZx738Nzvl6CD
EivYGUP5R7tLb/ajrHAu+2REbjj5jxIEwDgxwddUWR9Zr9S2Er0t1GEYWLyMQnL5jXB3gpruNr20
xSIgGwxPn549H/gPzhAxjDSH4VhmDKvAxu0xHolb6TkAgXZJFD9jNofoFaqMZkxdnBnsIH89SRiK
JpPDlhf8xTuhESDrGToTieY6zQ5PjcDSs+6FoVp7Ys+HUWmWke3zH5molidTAzaZsJEN1dXokbne
EkpECqSa+lX4O3jsPEnBO6rUy5EUmNHGdmvfKMcrlgVHnYV2cwVkhJYbqKevX3uROI+jgMUKo/GD
FFHjwXbXFs/t49vJboQnBQ2TFWgv+QNbmDEUIjsHuGaBsY3261b9Cx651v5UIrZKUn6zTCBTrn5u
Kv2uo0xJp7rYDG5V1Hya2IUPfanqnWOSHRMo03HxvgTW2QAoRdTLOQzEpJtzg/i4RkpoXLA83WFr
voOSfpTHYuwKomEVJ1uvygOaXMwmdlHgXsAd7F26+OTNmQ/LVmazUcqXSJNKCUlQGdNubXa0USEe
7DtNlqwO7gw1a7SbzaXfc3xbfKD8pKBXOMsKMCK2YYrRiX0ez+99cYDjZOZcx0r+DajmK/Qofb84
W5JCo+0oAdoPUPadvPS3Z1nAKmvo67IejKZVZ6Tjb66/7Gkg6okY2115Qf1HYqxYG/jw8a761Owm
medRo1LQ52r/NEFi5NAhdcR2bIRquzS5z49193dj2q4KoGCR5I4crBJlY8IG2lHlCEL1+7OZFgUV
6y3S7fNnPOMGMjZwdKBrVWuxXctNCh65/mnrtjAfTgWxji/7ZGkS8vNMglx92MGS24+NdOX10A04
0yDk2NxqhDwqdX0qvYGb2pZYnEt+qQ2wuKgV/Ff2ZM2f9etUY7ysF8e6lwMz4XrYR2jHI4mA86ot
34xd1a8E3ar/N6jfuMBIJipJfhxy5t2PV4SC6iA0mMouPxbpe+qvjbTevYIO3I8lgl/eCAH9W/+T
W04AaGUeZRxIBltrcw3mHRwmTNSOxFrBDTCiXiN10Kau+MrNqbDzp/08FtGtzVIlolMemqN9kZAq
XGPkqG8AqHdGt0klkuFTrytxZAdjpOXjH8nvQuweW/RwKIeUPsu7RTV4NzlAKYpxOY5B1cJwkMML
+HNuO5crpMePWAnNpIKy+ZhQitCkNBllUs7m2WDHsyB3/DWku4S/8oFbGGWj1tStMvDq0vQvm60/
R0Q1lbckl+u8lA3UCXu2CPKro3ySpSkyliyG4z/MN9viEixsyr7/4TKK2A+ulrnBKWmpvPzsN50/
xSjL0VOEFS9AVXWitHOE6DWys0yya+XpLKa40rzqDk4F2zaA1cCE50lKO3mvDQBmhOq4NUmakoVa
8FRiPyTtqugaIlYlM8+bwNM0H9G5UXcaT6MHvtQv+j9KgN39K0ZLiwBQgYLmsg9BXjTvOwoc7fQh
WEGNpyX25EqnL8Gg2VDzNqaHL1nueemdSP3q19ObOmReC4MbGY4w9dSgWGe6MRGZwPGk5+nyiIfb
8cSYPyqdzVgGT94pyBqPUqITm2VKbHDIcRVm4jWAo61DtEC3z2SfdBvDmUpi2q5Tzr2mbDbq/YWI
zOuuPbm/eom/EYqmiNAWWwya95ZNI07Ryxso/ndNJSiattbc+ysd+5U5D5HE0HA/yRALGgoTCCSb
3/8bk09cia+ramA6VRbNVqpTEY7lheEd1ecYclonmygfZSjyP39HjbBNC1NbOzUJbu/wm9YYJ449
YraelQp3XR5M6x9nNFQE6LzxuFsYAyfSK8Oxn6hKgHGVa4CTGMrThfpIFtxMnBGoqq4RdlXAsGnO
Cx+tD1Ol3CSw0g5cPrqY3Z/kEArJtlwVDmHaGH8nNFJvf3ocbByB56OPK3qUCYySyRkN58LfVYBf
moMzZ8/cPmlKx1Yhqf1sjfNt6+1MSwTPhgBrMgAIC64Xl1oCxcro/zFjeZz5/cAgOL0/sGcRx+R2
asieckNjDV1MOeq7L4r4RICVZ2tsCiTqJWrWPd4Q5z1bJXERWcBiFTQTkneIOOw0fE7wt3u66mo8
5PvgpqzOg8LqWdqa+ONvUgG0ZVrN8Ixb5htGDaUuxgwoQMh3Y/5dObBd1e7Oy11G+rYuJ+Rmzxl/
xd8aoFIV7ePhq6vf+ZyD39LZIEvYTdXPfZK4aiN1YC2ndIjVcBKv2rkAuNFM80lofVRgvUkQ4aa/
ZJJ0HyVbT0bTRaIIcAinQ9R6umUxrDW5qcEjAB3fyYet07In+fjM4uMRF/ZMRiiYdbw4cOPU2HNm
3DOKDJeLQgHKz21yxOysPHR87kc52HXTCecilwKrxvR8VetNkOxO+L5PBjjGYv4FubA5nxFJRd8K
4MuUMWIFHr7cOMuXd2RNGiaJAg0B/sCHQq3dof7nMtQOfEvfwaOanCox7FJdTSkeq+Vm5YEauuNA
LhoDdvxUuK6BDVWP9OhPss66v5D75H0+e9W8mIoicDOdHUN8h+MGy7SgRA6hGYoXWf7EXKM6Wxt9
7T74B6rAmVWQ7g5Moe2LOBqucMGurHHngD+MIFA3x0Lf5WZQEE8FffA+x9J28QbmsSYKuLYPZB+B
/YjHMO5m9zXSHQ/mrNUxPo0pM8cVpkJdYUHY/2jzHroxKXJysumyzosmV2XM68FMIPmppjUK+/Yc
UCY3/7jU5QW4LscInp25G+CbhfMkxdR0GROtF524oevdSe8bYFciMFoct/eHWwOnP0h2hDzKXBzi
iz/mPRAdNZoG0i/Xg8gJlGMNTFYDHvpD9dmwtc3UKyTFXEVr3aSNkugSuM98KHiy/bdUP9ytVsHX
bZO6JmbopN8IrguBQbBTttS8iN8SY0WzTpHgS/j2qHEL8BujGkQo96BD+8TeuWKueWoOa2TrIsbg
w4mXmGAvgDi+aax1t0dY7RDTDpN50Xox5aWavyYdsQMMF7DeT6n5MkEZDh2m4fl+qCrdvSQ7fD3K
fptnSkN61r1wiKrxCrNg3W8y6SuA0iRmu+VKFS8gluhMF5youXNpqs8V16tRCty3BsFcIPcS87Eu
2YcwkvG52I1BRJt51Zme3GXYz43BWbupYXMs9BuROvrmM46SQKEpIr3EI3rGgt/MIR0tpGixvLN2
ujIqOp5YzuNsNrtn14cOxgOkYuCcrhJrrYDugYWMsQmv3mzD/ssb1MDo8d7APLN4RnIvvPndlZeq
qrE6M2mKFZVJm8TqhZsAUgT3960JyTrY9pcGiOVH9cvLq8vyUL6+XtOhB0n1ktGD+lI2aw5Lqg2J
n/4bSPiSlpJQIU0U2cx4/dkI6zwNemS1ePPmtydL839bqmUPYtQZM76XyC0SPiQPvD+4YGeY6r79
To8E3OuRnu9amgRLiDBRr0gbPIHgSTz2U5Cs56CJXyB0UbNxmo45TifMRmQEwfUPfEZCFU1OUJht
DFvRnvqXPQsQ7cc9TIDbvguN42sntWdqBhx6ThbOOgVICFF9ZiYAaeoGtY79EdIIMSMu32PlO1GU
cAMUO7nsxQ4YUmgGiOCs3Pa2tb5A9kP3EGLAJH6+or/k3mXndyTk43kU1OJmFoFpZRZs2veYu+VC
p8WnK+pKTiMOYNi8bLPYQObOiz0YLdiQTQ9MX0La6PLDv6+KqDtt/VopxEsidIX88hVNMqEV3Z9F
+gepb3lTO/ppkWOhp1jkpJQs2SUsdguXHpd3JP7H1KAPnEvKDX2SQ3O9vGKNUE3PHZhq1/cvHYwT
ORZxSKZfZwB0UOiQaDznyBnHtI0XDT1N3GGlD+ABM/4Tto33zhzV+M4leQKR9gtPQzSv7a4Q8pm+
mNGrUwRWz74GE5Uanr0uI2/D8/Kdcay3awU9YZaSZx4EZZV4h9YeZ/r/XUo6cAV0djp5dj3KhPUs
91EgS8LpGu4D8ivs89HsxtYaCioPCr9mKZFx0bsRKEK78Vobqy2b2lrzZvDvR3uThXgZxEhKjsQC
TsGLFw/YCUg4C2Osx4WTkmTOFpZttaHznpX3eQ+4EYs9+WQvlRuftYDepYMSRULJbbcV5FZ6Jdc9
3S2vOv4XFWY4XbzqzIe2NoCqwET+6OiZjqoWADym6ZM0f0fTZbbsOlgGg6RB1uThhv4epnfbjKzZ
uCkugJfahOlywo2XDUzcA9HN0KADdHUujpIwCEM7qEjnwZcJ6w5BFyz6oEXayNng6cnzLHog7iO9
ppzWIgFZBS6RqikEr3KIhLW6DTdJsVS/PsF4X+qeEWyscKqaLROAsIBmrB4qRPBN5GeyM2cTIBIa
IkZRro802AXgnXS6Vx1XVkRRUablD/4RnvcDMV6H5AHspIvQlU1jAFiMNA9a5ZI9Z7zeRLXKKA/U
X1l0/eJRqE8Pzgi2EB8DoMiJ+Aok3t1hg2emUlVQvxcz8t3Tp0aVGbOakSxNTAjEiMqi55Q8/fy+
/pSvBm41dPoLDUHd1WjVGXPCS8HZBsHhMvVnxgpwVgoILY1Z9Qk7j0WZjTQvBJAp7ft5UjgM75pD
DGAnL0vCE6vOWS6Y8nAxS7FV81h51blAIj4oSDD6rdCvr4e7RbFP0bso9H0q+i1aKenECWHl3Hrp
sVFFYjbddVRaTdNszmE/1ClzPQhEC8ltNj3Sf61OxpiXarfsy5HslEhWjzalt3Ks+1hx1kfJhIE/
wC7pjLiVvJHXMOqtIxgIQhRGi+p3zsxRe/4LDR2pmhtgEg86wV+Pvdsa5dYrrniVr737+AemKMor
9mFU0VKx2Df+rVrICFW8s9KfQog4vlCdf2QhWv1qLPQF1Act+zOPxF9PsGZqlL+F665YzYFQJHyq
I5K/4yX5AiuCJC/JTLow6llbAGjz/9sgk05qvTWMPbIlZqGfFUMcdH4zaMygkVAHTmBuB3Yniy/u
SNoWKq/mUhWLvUQH8is5to/1MASe8cCYMdxc1SAqcSjjWI4M4uy8Cv9DJWUlIQNDLdl16+ATVap5
9X2L5mQ5zyjaJCDE0qD6f2cybTURKl5BGLaqIbmP4USKzE15dajRUqnx0R404q/QbY7Y3tipQS3c
XyerQe3F11seKqKqBxIZTJuPhbjWnPjb8QgmrF7bXiCri00exoQ9XrYXYo5WejQUzuGt1YhSqUu7
JgQP0y1mCdTgjn+mZX9wlUTVFKOZp6M27RWWYeu/I1CzIyH3OLGfoIfuHwV5jaMfm4NxW5jy6YSA
BylgaxrIQ/Nkfu+4fM+8YBrvZOu81rs+24vMj4IaMR/wC20JT6YWuTOm7RSjxTA9Gre2LuUFm05j
brOhHXs8+j/1f8pPW+BuoKtMs559/F77FbZzeCZv5a+sYsa37rdijTDkm5V6pCFl/dSswnegAUny
dzLl2RCui1XdJ7hdAuTJFZmfweoS5FJLxWh5q0QJ6pqeUcKNMZX3GHYo1OX2nEPBJn5/CUDSIVly
Iw6BbAG960aJ1yTCr7jZELPnaVnZbuk6+Ms1EqG5ULaRv4G1EM3VCKp/eklXHlfVOO11DjD61lCo
QCiI5jGJeo9tfLJS+OSOVnrKjGtjclse9kYbhwStrdngAu0DYbyN9oT/3kCzP3fqIMQm3wAzWeim
8I0c0mQcJfzn5KjlWgzTKbI9hYqsqNXYYWQ57/hpofw1x4H8gRonAbafCf8WK5GH5S+36cUNd+DN
Zm//VqKHL+NRcxCjGEI6EiTtxnRGbvncS89sCjxtvz7MQYZfDpyMxj4M0jlvvluOHnY5rBgpGa81
XFMSOtB3V9sXil7QTmE8yz4/VODMVXEImbsT4NDJXeXVHMnTuHv/4/axmnoozolifWfZ0+IBsWdA
65uq1R759cTUSctqGV1L1jkS9XVL38vwHbMwOrNBsbArGI8IPEUJy/jJ1DLmNNuAXw+3y5hsf7jC
I2d+BeVSL74f9fqBByT1gq+X8smgpb0wydLG4AQhR2opBqurOE+6rYg9Dweu/vtKGWtj2Av0sXT5
46dq2loQUsvYTeO0ZauJSIN+PnHPGrZz6WKi8u2clkeVZx0jSZzbyLwImgVGi1wJ7VojwhlDYr7N
OUB9qb1LxV7au+03SQfUBiMdjG0BaIpeBTRp3TxhcD8rwH37lZRyYFX5sEa9E/ZsXym9Pi64hy+E
JvPpPLI5Ak0E0k/03q58Y61fZkaclqss3XpsgFM2yGNkZXV/LkodapqJfXZp6f59Vqs4tU79qjSs
EJ3oOJVOkbF8mbIRUGxfK79lrLwdw1qdTPhbAxusEursUxCUrGxkCeNKtggjWkl6qJkX3up7DJ/4
5sUqvB78VOHnjsToow1rGtaqn4yO1VWJyWH6/hE/ao+Axww0p+oUnIfjsNLcYbA7bAPi1Hnpm2ii
GuWtrQU5CSCQSemYmVF6TT9F7tqtqQ9JYQpMf5uh6PDYJBznpQk1Z2UP9ySUiKQUtdwL439oy2Zz
NUKWGjaWle5LnTiLyt3ImbETA1rHzb/ar57f+r4Wz0/htfWq4ZTvQpjkGwP9BrDG+R6djnOo6Liy
D2DX6ccg08X0AE3/ijSeQU0qzTMPNDwCIz4AGJt92uhb2RTw9rcche/qZZeDTRkW6dJ8KhpmLUeg
JiV2L2uI7IVsQunPLjdDkZoRdkiesfNVLapdpjgc8jU1j4dVr9NlmN8CydBOFsiUKmIgh/tpbPkT
t1J+Takb9VDBkXxEzUzGgcZSrQq+bBbUgzpa/1aCO/5alTN4vpTQJgHXfWy5ToegqlOsIfRcnBBU
5lNbpgnoOjZs6k5ThlS7xdvCONjYS55bq8ee4nQcpp/Z6rcQoFFcM3ZQIv0fkKiMmtPcQpj+Dtg4
uV/at9u1wSRrRpOO3x3FfdyN7jQPSeatzJja1/SF3nEUkrTu0iiiaqiYF7TMcubB2O8662ugaTHI
usGSioZ/fyYeCydZSXP6+WO/s4lP9C8ZUww39q3JZ5TssYZbFQayG34/PgI6P44sD4AQEc+Q4z/g
T9Jbhs7A8ThQuevLd76VJTu8LcUt99jZt2YzWQZAMihN6tOsu5MgrIvo9ym6zx6fhAkkAPj7fG+m
RytgnTRk8WZLWaJJly/hGzHed5hadzfGlK8Uy2jbD6sQEVZycaeBTqhpYq9GlYrntWcEnGji7ttj
iHhApxjI/wieNM0EMODuFj51WkDl4gtd/3Yn7R1ALMsCJjhl/YtSqXxT7hT2RRjUErDuzylflXiu
5XtCOWOK1LW9or34bVg58zrgP9UzytbRs4p74TiIJ/kCzvVwk+DCaCqWpX43K/8p+pNGzJTbfrOz
RvFRn09RnfujDQMjjWwu7GNfnKXkjcx+mkNK2CEV/eZ8fsvLQLcnvA87LQXRwRfxKm3I6tqqoEEq
p+TocKQaTlii6SEmbJwKd+qE4M8ZLS8dWYjtfunBt1/LOc7/R6htt18NnljkExoM3fQ/3IPOrvbG
Mt1TuZxIaOsLhGZ3a3weRfHftN0P6ZTLdH/lwCGdiX+DdTJ5hqXK/glIMb9CXJEcMaoh4v6D9/ST
dmcdsa3W9l4tNMgq0lR7PPI6KjAe6LU5HFLeW2ljeYLfJMlOolYDYmg2LVQ3mPQjhlQj2u9/kDon
UZumxPEXuXmxjBaC6sXIAZh8aN9y6XFuz0dtsiTqC9rbHPQOQTt/RGJS/ZRc+W0YoBg72obfyBQv
PpYgs63rFGJu3sO7lqDWefnLYaAiyoRq08J+eeYC8ifyOIT4zZn7jxW+fIUWCSAoOOwCtPNe1Luy
CWwB5btXe9Ihp9SjlHvBNbKtrKEeaTrliRZ4D9YEraUrA3/O+ZrEzPgvtwb7NMqbUmbYOclAHA2F
mMMKhdeS2oE9kP5qdr8MnZqjK0sHz3HpiMKIDL7LPjkgLpaEinh0EPRhqWjJpSMYAxAv+OooyIRg
+Bv8GlnUyoVvMOnvvoApc555pafIbvxs2CUmPfiwihEN1nDlk9CL3x9Bq2F3VDLsJOGZXuVNE7Ht
v0ubg3nnRqU+A64ldYML1/pQROcEsLEULMqVa23rX1Eb1PtJ6J+1qWnI1nE/oimnScO3MHfNhZfw
J+cWHPJTUMGFOItvh4QQXeinH4sYCrvNucZQ9NcHV6kQiOKGbBwkDv65IBi/BrqlR80tPdDl0e5E
gMd4gtjbVgV99QFEtrU5hxnF+oGsmANHubxwK/FqKPgNgKH7Vi1o59BnX40gxTtv88GZv7j3sAc3
Xpqi64TRgF7vk5oddSHQwa222V70qwZR+alDb4C8feO0giXaoKcPECbutFTDcreMQQaszE85YxyP
gKP69axAHtkgMexuGB6pZNIDl0OEu8f7nI6yU5+7kQ0Os68lE5bbbWI/jF3x/LGhMpw0o0GcVPol
mmyOy4PshXcYDOdAiKO5mdwUJkD2ohSKGnmJibdO6tBK2r+cc7wqt+/38+zo6L6ixvgtijUmpJuw
7VWYx78ta9eCuIGZpB81S63FGIN5IVWYiRYNKY8Abh6+32aBorPhVWilVLfvnbtf5Vtokzb4y3gQ
rBcq/Rwe5oVnL4xt4714kVg3FMB6j/k64kCLYkCvKZWDR/HRGRd9bxhDKKX2SjsmSsEIJ9vL/4vd
eQwRCJkl81b+3VQHscGtflIdGy8AnKQH2q32qc24Rc4HsOTnlJ/LgpJBI3rBGAEZE2cSb5oeQskk
Mz9YDZLvEcSb1Wb20fGR0HAuuo4Q5Fc8jBg5BuWWvDognjfckQMfKHqHHgRab8QeFpMqmFRGjriZ
YeGVCU1k4TCvV02jxlJqaJ73TARbhvAS8aiV5ucnbArULBzIA4tnJ/WrFNe+NpXATy6RrKSadUtg
HpEDDNjlkjZoX3UcAhIDTQjdy/v2e98lcGJxViYM2KAll9Ep/PYUUox7C3X6nEHNErxh642VylSM
iowKosFhPXtU9wYXeefMLSv40m56bNF4KYXVO4sNyX6G3W7yv3D3eNZcon3fK+nv9hfqR7DD+5oG
gVPetIKDktvMX3W46vxDxryq39jZiOPxM9iEtJNaIOpkfN07fLsnoR34uzDPQ2M+pn8bJGmEdqlP
0tkX+d3/5OvXYeh04xGTP0t90SB9wT0kaVhiFM6rbS52eT+QmBITbObhnAsTzJAC3ikqLuijqsF1
BqsGKaq1q0fTgNIqq9hvMHlQMrpX3EEqCYaGYskS1RvW/AVzqyqLhp0FzxgY2IF2BgclHV8MO6Tk
JOIl40GStEw77jmFkye6hIwgZM8pQErs/H5Tq/Su3NtHiyKn0MrwibxY9yjEzSx3ZcJFZQ49KVJF
VgfiqXmro/AwZzPtlIkGP4mmTXlMj8+LYdXWRr4Ix3DHR0qKFJZWrI87WY7fb/smn0uifla5YF5e
LCupXsMdgZTBa7s5HRbsXpQIxOda5XAiRnB3mDq3k/fZsYz3WqDJzWwD92KrU3fg4PhNHQFXrWwn
LzcU/Kz0byAOq2i3tXQ7eylAv42pJLQJRF5jJ09i0fKvYCwz2sbJ81WnnVeVnMXJtSrKTu/GtXvn
goG1pHn/Ux7kVNqMH+Qy5nSq6Y768HUdxouZ//VG7LgSVFJaiZwrt+KCY+pq90aOK1GRU7xEJOMO
ZLcQ2mgWmKWmSnZBYBrK9epL3Z9wNXFnp3x0/ber1/r7sCmezFqU++hXcmyeSf9mdRu0g+SKrYhw
UU7owmU5odS1RhC4rWTq/hyodLYHpn4tp9V7BcN0fCRzhCxY9CaiofJO9c2Nu/xoEsih1Bnm0VcG
SnM5vPWUQYx2bUR+P3+2yalpMruQQjRUPhwgeOF+Z4GEfuurJAHh6am2KSxQZ7S1QqInk8+lWoTB
GCaEq5G8Y0pqC6T+QC+sDquFoHlrLFCJscCJCf0pqTCgG8F7+UqmGncCzaWu+SS4Cbop/Gg0/CFq
jWqTCCmy9i2WeZGp8ZcSyp20zN5+1BsM85YIv69sH8U0/rjBgIUIHtvoFJQz0+qVU2sV7T7kJ7WM
exSJMqtSfVJRsO5GZFxlq5Ws7NYNsbhxKNSYw6tqHXRKWCqVF4FgB42SSY183iiRLti2KfRAi/Se
t6bzGTV8HptSGzVH91xuBU9KQb4y3D1owF8wyBizLcvllunAdxpK0tS7dlhE86LtXKg1i8/AxN9z
KdP+eXG8/3CPna+NfBkM4Et4qggKuNN7AHh+SrMgMqofERTNp1ZzFXvlU+KDcsG07Dsrkc9kjJMS
DqNIymrrOjjv6pzutsp5uFsl7BoJhhePw+A956GsHquXISTqpFZLPKcGypNda4QX7Q2KCB1sujwN
2Iywr2J0B2uO9eoOmkrUGouj2OpTO07vVx3517FuiyBn9kZ7bpRpDKlAqm0IaZB8y9KUsrNQH1fX
hsYCSsT8Npf2/irhuP8P+5CJcMnDXivEUkV/zZJng6vze4ih6tpcdu59hSZeQ62fGsLxioZiVu+q
xt1u7Cvctz2BGTrACTkvZutNC2dpShwTtO6Xd6uj4kNs6uUvxiemp2mY5g7ktsxoi8uwXi/J8Alb
LViWgxJ17WKEcFuz227Znywn0YM+Y4Pus3vSe4/27twqj9S2beGl3+mf020JDJDSgytFWAmLsrST
/PBRnJLbE/CqqOh0YlQVuvsEqx8LnEfPYfWBkm+loTxeSlS59DgC/vDLKNiyvUfSMLp8ct8pXZIJ
kWNKvT8cRwp71z+G6qAlVyR0YSHJVqD5gEoUT7qPXNnXfXZw/b7vWihoZA18cePiBsQVjh6gHH4G
Mg4us3CMh65tXYYaq1bLEV2RLFKvVeZCn7uiOBPEB2tKtULbFAXnWFRCAhHgwfcfPGTkxGM+JPUY
7I0lswlQAXIuJIWKIkIsr88q2WaNR39sisARLwC2YCxrM6sRYP3o8crpYlazT11Bj/Df8XrFjXNJ
fCiu/S6MdrSBTj6BiL/mIsvDvN2IUvmSB4VTS0HMungSUOTZQd0znkiMDLouJx+/rxLzOPLTbqrS
YuRglMFryMiB2Iz5RKoWWGtOpdOYjOhyvE3l2Qlu9ZN/ULPk5EqKU9gNo/mp2Fm/juSaNeREZRuC
pfqxhWwXxQ+mi8vBjxb9YE9uL0DC9JQe2ePDUCXpQ1jGMUBTjQFTbz5patzVkmTlHJaVS1nDfXfK
Nhoqk4w5sKmjC/ZyOUWHq5MsvL04JO4dMkYdzVQ77n21G+ajkEns39FNSvI2XwPZlcsGf3T02PDF
5nwiVppl9EI3o/6Go2u5p/nW/cgpRy3oqLw74LJsWpIbtYhfW9XdW0wHSZZDE+1xqMsD+bsSWT1n
aRDI45uNkIkd5Ay7zxZUjJOcJAMhqhsm8QumCZ8yqBcDWD0mmuEIVZZwcq/qxbMxeXCp9l5XfVbF
A3D/+enRCa/8RhA5N/Hwma5BgwLkYA1BhtZp9nwYULZVpyrwKeugW6zRnjMg++UU692pIzunkZ2W
Dtr4D3i8plC5eonp1bwfAUqO1KTLmqGJ6pdRrMLRaXdfrTYrOIlU/D/grWaNAE1JZzx48Mub6kaV
m5526L40ibSyEU1eKzq0lYY4g5/Xx7jHAbiAZAAj0M/tRpZHO4q3Pa0xNozXx3A3UsNdK2IA2Jkq
Qt5qYtfxgLnfwm+UopAigBs3tKFHQNylDp1+0e4Jg+DBg+xfcblP6oOu7GG5ZPAkL2522vkAjVWW
lVzbihSzIuceaG5ebjQG2W20cuLdq3Yl1jsH6syKJRdzYSFAMd2vA7FXT+oosObE6ZV4y1pBkMTa
wnq0CMbkjVUEumU7xnb91NLVW07EGzQUDn7ouNXnFSelD24KHRFsyH2D9EVx5kvhSrc1e01AgBOX
xqibwflZ8OadTUH6zQskSHgmi0Kg/BUiVyEjfMHiGwoiR722oxSiWNapccVGMgQKjyu6ETgZr1Vo
ebkdbZNFISrTwiotZ8TCKlelY6e4z9pAdxo7J2d9H0SWNCm/T0I0zlUhaA/PcF/4rsVXhAdozot5
pDT1pxTOKdHrMYYP7T4s1ZdzHmXKmtA9QsQ+w3Mrm0rGE4xIUxBp/fulnsLUMZrmAp7Z/hELEr2Q
6qe/LWiEdIyUjln95569BLbYC4Z4kK2eOy2yKd+9ffv6M6DHkKyQHAOAvAJgwqeuYaOCWui9jIZQ
K55ILosn0onVFwVDoPz0eUNcF41sbfxQNH6v4FXfwIyGPKAdmueQ04xGWj5a0esK7SQk6RG9VER4
BwrTFNOu7xes9OhkUwfst/KU/EzfrsaNsKz/ynhm+fzQYveSy2GjG4BhVj17ySyM9jrILky8vUaS
j6qHjZHuLu03yXu8TVwd/FSg/60G65hxOPuwmze1kzaEcgWtrX9AUf5KxEN1UOSVbUcBR8Pakimg
Of2xVH7WlkBu1fVc7tX6dVOqJdwrrouT31PqhCMet16lAbjod0AUMIPpEjCbIAKpzbvkUmJNUspF
kxql7dhYYVNZ09YMds3KrR/XnQ0V+kZlDQ5WpkvUo19pb9+E+Vkn/yMobGznnu43bMrtLRrGaH8j
zeE5rjddbLeCpEBlzbuOoVoTc16+KeJC+76DKE2QDRkqY5aWtp1AfyI0LLNsxZEfN/prWpSkbGqQ
tyTXatNbom21K2lftUXz9rjjTeKB8OT+nJ1p4vV61T4hOjdNHpjBkt0NJCJMeOmOv1tqdN83YYbx
7fVwXzJoPQ2ONXPMoKu/a3TiSqsuz0M1vT5yZBBV7WVqq9UA+5ZrJp5beoGwyU8FOKh8756IFjp1
hvhfVeHlUSa1mg5ihJ6tjg3E4VjlsARNn33ZOXgakn2PkeM67TSebJoLC8pOSMaS6GvYc3iAOyva
vYoxYn329dnVJYrmNy009IeOwrhb0tUogVR+8pDyO97hjBH+gnNSM0/stWSj41K61Fw6xHoiNny1
TP67vTxMXkD5MqGuCJJT48LzlYzzHrDIpNTfimDYPnNXVTu6EBqkKL4wYM+FMORxs3DkD18tEvZw
dtIkUv5iQjKJ1wGDnylRDeKkY8zyME8GCNcPQxgm/JH0SisX9a2woiIXyJMV5yYkKxJdmPy1AA+5
OTxh6EU33IpmG72qx9K4w3G28mH0WbfP2hZZq5WmW6vXMb9nWBdCuoaXvBORGi5bVCb5jzYVtpjp
ftfQn4GhG6hoDxeWEDCgGhMiDW7nQAJAORuTmNJNNOc2IL0/Gl1wJGHt+3/36dOJLupAOlGKf73o
2QvScwYjgcCBYrCw+kktxHbxzsbGsMpdAhH6sHLXaYBiflnF4NFNbRLvxQANij2b3ivtyZ22WmRD
LaiSaqO/nCSn49jKxEviyDLKvPH2JCPGexJhkAd/VN10FJwGJW7x2Ms10BvXJQ5drHOtS1F8FHH3
9JkQ/RzUdJLG1tJQIGNU0P1v08AfnkpyL5T8p9Ci07QLFS8iqnoyvqccLWckrtWrxsu6pVsCtLvU
7+sMM+X9X6JbxGTzH3H43qtjcQ9R6cnUVeShJJG9yuNiyeOVqvEAf4RNji0hHNtIxF5WsXigAKyf
3I6IR8zw9eI2kfhisOFunKJM2V2ksX9TOT4s4wKWD0TYWTdv9yeC1uhIWSNlaePdv1bLkfc96oJ7
fjX+eVHAhjjSLx8JEyRzQN4uCWz6sdN1noo4oqIGJGnU/QFC7vXvhqPaCmxePKCKLM3PwdgT2Py+
WDPQJum9wkoXEf7zX6rieLy2PDAVF8w/3bjnh4DgNH+P3iH73rc0d1gw3gvD9x+Btjq0RGWd1Qbi
98X8xRY0BBYI7wOIKkZZyrJhLaBNBvh+sV813UkCy4hLqP+rvkTDM4Oi/RI3lg7zeqvvXR6d4Vdh
8LRDITdd/T+4x9sgf/qRf9X5W5/7+t8/X8bPO4s93JALcMx9MBP9kcQ1Oi4EtrZje3oWzge2C09Q
QkRfXzBNAiDH+T58n2lecpSbwp+yT50QX+T4Ezl73wdqQlPqotzECTLMwBE/e9xDCld2Jf5vEtSx
hjTpokUMVj5AZnMLKnpQ/Il7zRZjRbj1IDwsTw0cFW5I8WA/ELsLHoaKBIyqZaNi4+i0GvNLjs/i
wlVHtbSmRQSF4h9/mNo9FEbh1szj+lWhDJ8WBRYUGq9s13e6WcTVAEv3lp1hRDFx+p8vLnrRDBaZ
el5I9bldafyHdhFDi7PECAgO6ZZ+Sb771up9yxi6AMToH2QzwKmV6bGwQoaJnx3sihm0WEmxuiuv
qVbvDpuyyFYGS+ISNolYMfBLTrC+H4EcddVZGaun1FppARhig2L1OBANuTWR266Im05JMiBnOJhC
1WC0RiaBDzIhrL8bbxOuRQudD7YIutRUGggd/ZQ3D+oy4jY6VicxdTw03FDPYQ2OJzAhAej3LvGb
CCwIWvaIknmyJNBEEyQTkSwrPv9VAdiKZTSwOTFR+N9RrMRUkXje9s5YJ4zvCZkUaX3l5HAqKNTI
RDo+fHN3y1DgfmSvLqLY0OmHjeU7bQezMQ8fMb/eIMxPxSCMYtaAKkXtc5fPBXzzIIWgbB1sO7P/
MbGyl8ogDH0QbtwNqUnDbkApeqU+FtIf3/ill9N8lOziw1ibTjCieYeDJWXkB1kSQ/ymwNG9bO1/
PfcWJSWPSz/0AOmbXxMGbcGZ/30NxPBCdKwZZ7lajAlaaKqiqnpuIIwRsuX6APSOjQSCZx5g8FR7
VAC+1VrBm56+GgZl6oyHuk5vLMgSLowy2gCfFY0nK68P+uTVQZW2bv6qNOdabQOMePBJWj2uY2mI
Cf6UXvmL/hWLtznfbrQ3YnENcXFo3euMPdpH0XCEKv7R+bTy40puF5eBT8F3YDJdrEz4immyNFCJ
UXJOxgfyH2PV2Y4wV58UAZEgcmFhzgBlsnGCjbZu/YL6IEOBRqOABz+lGQoFFuW/9PnrqwFBIFUC
IUy8lIQzGlZPbAK1Ykf5p3L+x2ksfNwcfxvhEDMc6Wvp0KSJx17pAnR6Th5lpVDtPvLmfykBM5Kv
RJ0rtHA12b8RvW1K7JwdOrIDGho4Fm0imOpi6f2HflxUHkfRRSCAbRJY3DcAZpFbjsrdhxA8m8CB
n9S52RVFTDWsrG0qc6WT7lpNSpsSYNFP3WGNiBHXVSw+0WvA9vFEqjSed53Jz7zK/kTILX5TiofJ
pSnIgugp1r9T/ojcA7f6syDScZyNC+PedQuFIGRwabD7Eb2m/lb8D+STteGOmyxW22s5R6URFfXz
EmwqaHXMbMzEkx5WD4O55FBPcKJuV8jT6ptEilaKGTDj7iPaC91hMLdA0GR0g/XlbXjTCT9ckIFD
Zy0SZlE3XWatgTw2eYyZcZN+5r+JrDbHYF25vzYxTOkynJ7e/VpowTooOS5iSjpSnt4TB+zBNDNO
df1/LanPGC+7Yx0k/O5sy5TGtCXrtqgbcpo9NFXSkK7M6GRBhVdPxe8CxVQTRCj3KPhsZ1xSXb4Q
deQelH7JV3dgDzUJvoE2FVcZ8gVhXyMWWEGVq/i8aHyNmHDDadjIaCCC3bPO4K6aOtzfgIVo5vnh
cx8fFOhcRoYHLAsrsqfI0U324ND7VXzTHi1PJrOxqOzAlcFZoFvEomkjuFlpfTJ5oIsTokTmPt/Y
JEGFu2BBY7wnFIMfxB+++9DJ1v3mSRnfD/trzoLqpNSQ7G/RUYUNjEyqZR8hd39NH5WzzwRDTPi+
Axgiz7VZgpV8EQbZevKwE4hjq6nTCBwIN+DJNGE0iuhSWuK+ip/FUtJkbqImZ1WRhoGRVq77ToNN
EpXHYYaw7weyNaalrlkRLk76HC9CcMivCi44DJQX7C6y9Fu+/WofQeNyQEt2vXFFh1+7KU3uhERB
C8m9MyqLYTFRj0YqbunNRrS5lnBZUDoX5FctrBd9UUCmZVJe9k+KD/a3qRpjHUjIsreM++2KeU79
MmkZTilyn7hLnBLNX2hQVj/O8VfEaOVDvWkpe9LVShZU7G8ALUk3PEi0rNxriiQXZFatZItssAZq
MBSCAqu2YKhRd4VmTfc07ysadM6OBdtxOjkjItvh+b407AtmgE79WFK7I1gRpadb7UnGbzmzogpe
NXmYSGrT3E6iqEidMBQaaG+Qza+p4BZoexAvpXes/O2cx+4ZV7dSxD/oB2lPYxwPI6fUBXW+ikhi
1hr8z+oHSOevmeYAd+kulelUfBrh/6KSqnYCJfFIwI0AXcQuJqKQfMSzJDgH4+psHaoth2CsiaNT
nSdnat+2GCvhWfomMwLKna8XeKOYx2ycQhKCsLIDT+KIzf1HoYQDCTjQnxW+wT0qa5SkVYwjeSO2
sVdeCuHcDkiTeUqJ/LPR9f73zZBN1nDInvDCJ8GaSQ+uGvYMSWl0yDNXPPl10IyUWyNBsmoiu5xU
q0Eo6AUCXv8V4eMXIlTRbwEiNJlJISygMHlU0xRw4z1seuUV9ezdFgkzLcC/N+WQybtIcnB1ZvMm
YYTwKDNtc8JCRLWEOA5Pb8dRDht4XvMmkK7fXA+cC3ZMKRVCHjR8BmfiOpfNctO/qMLS+kU9WmYJ
SAyn9t2CN7jXbfIC0BJEN56ALPKD8+9MBK8RzPx/ddJ/N6B3Dc/m0ApcGdyMDqiRB3p8NPhjhJnl
yUxsG2B0H+/1+HBw8wrTv4YwjJZ/NeH6ixy89SL6wZus7Gvd2fKiRIqDtNERKhBjHy+z+1zL4+Bi
AfI7FblRTKLcJe2Jm8YWCPEmDxOSZjJACg6l5wJsS51l5Hx5BQYEKJp+icHi2PFb3aKx1IrMwlGw
hX8Ji3w464HOjMBbNEPsVdl7MQJhGNPjPWdN4ffs3kRxc+NW4bqMfTkInhDhw4AlqaVmV5kDQksM
O/1ilqkSYsgRMeB96XPC17ZSpVl9AFkEK/3CtsdmTeYwz/EJUIlM+BgXmtj8MCP1NNNfHaldJrcH
q/zSl7yk7gNjO8yc6G1ihtqERdmLYwJ+sFfF7NuBV0+0iegAK0WpUCrwq6b2xbf3YwnRgAB/VQe+
QDRYVRTL9vHq9lz4z/U2kGoUzswX4j7hsRP766YQNf1dxG8RZSlGto507/hX7gVTbSVoAUK1zp9m
/pY1QJw9WDd/6sHKKGHmCMZpvmN1Zsbj+8oaK/CQxG56XWuNpzAbFiuZP09GlReTdSKsYcX1kMNw
5qQERPjghjVckNQJW1KKyXm01T0LEA+FtQYjPcRra6P8uMRYATDEPJCcQgxn6oNl9T4m932I4x6L
bbwApBPwEnIg8r7emSnqyvz+4SaSezlCqM2h0sphMRUxLuQhtWjKEER1A+T/qcmr8dEj2J+UeGpm
MpwfYrm3OpJftRktlugG0KORtTpAJzhxB4GJovDptCqxOl5hPy7VYhZzMkoc/D5oV+mBksuIllsq
SgOqbrz7RKR7G/TJTwLSH0f6WC6XAjmdfIrif6MXwZGe8BspcjksuZeZwcXZHM4rPWefOsrbkJZI
XtKBKOazR3Yz2XWRW+cQyGdD1mtz0w6lZAfUBaTOHVsVhlQ4TkkIvQsF5Zf0/SB91lU18bMt1tAs
0zpDMVoBv/pQaqkL8fGSi3LgerQrOOpNYll0i10B4st4AxZGxUAKTmrKQfry4g1gHZEsZoGSq2W2
To8m6+1qstskNClW0G+5Grn4t42mVpB4pkhxqV8Dh+vK8CnSORACmBPiI7BJCBcx+Dv7POnkbpXH
6W5vtrR2ju1sVTw8oYzSUCCiP41CTiESf0P3ohKM4cm44onfNyThQlazBiILQM1N3sV5VDU0RYch
eOXPAGas8g4HrbPx5jilkI2WG6fuzSBCqrb+ACA4NwA2ykcIF8+kwYA4Ri86uzmZFEm4QetGUgQH
IbBgdgtXf7DdAlJCfekGpkD1TJcj753j4jFWGZzNWo5qXeslDg8CcxAvh+LegJ2GV3XtokhvHn1a
CNN58gMSABHikuMQQ1CSyeiELqizLt4GQA0cI/I3TtGTJoh1O/mg9UnIygbn3UCgzSkxXzKaQU6M
ZzIuNkn25w83TY+M/XCGqFGOupuJj0hWaEKfXzc3lY1/kbAeXhlFUDyQl+TqkVZkQLhCb0GFlvUm
P15jfQxa+xrPcF2fhOjlg63ifi6/OPV26S6sycKaIFaBGfdPQhpYSFVkq+G5Krfls4Ni8LN9zvYU
HZimb+cUBsoI4yfHx1I/h+Eq7nbwD9i8iptFkAlZ1WjQYo2i7jgARQh2Da1j5Y0ArPT2uQzyiK/j
IiYPOI3Jos//Iw2vSAs40YKlppnoSXlpU1+AaArkNSfmlLZhYGOCksUSiCxFhO2IYKOWXAjeAMsL
QvfKrrTymz8LUda3GLBIHrFGhhXSTPTd8ltxrQyEy2hMGwH1diBwo62otSNJCv5mnxQUlACtHAlR
ZWvppv6DWq7JwsTHOJ8x/6UxS8E/lC9hTs0LF5bN2ssR/P2ghD+JAvAfHJmQtXF7Clp0B4MOoIWx
CHc6XsctxN7i3Guuw/hU4lAO9gw83YTM516HWME/IHEvc3iJM8+UYQXTFalN40VaBUdJ1o8og4lU
Pc9rh2c9+nncYljhwUmJeRkEuuH/u7gLxMSvbO1hgKZyarjqihp55M53b9+TmryTgfaO6pBRKiuQ
MuQJ5gn92U3PBvmEz0Qe+OOhr1jCu3oB4RATgcVJ8Du9+sReYsof036zPzgCmwEUVi+/Evo5t9Xm
9RMd3DvkAuE7T3PcRBw4wvbw5mFe0qBghC9PexV0kmqJPCVWsCBXUy8GYr74P3vB0iT3e/bFzzVv
Agf9SDgrSJZd0Wly7cJWCShgVzcMxNQ6mpAfh+MbHK7kOcsbd6UFeoFOL+9IDet4sKwZBWPh0EYQ
wAzmdSOQYOvS/phiRu/jYVWP89GTpOifKu3AHWQvwwC3/zi16ZD95orStE/ip68ouQ+79BBQgW0F
Ab8kM8ggPl50iO69V9sFPi9SG8S/Zet3qK/djDd+RnA7pHyZcQFTLcYfILJtdReH+xPHE2N8QbNN
m2psKbRc0a1uPYplWZTuMExTgZ8CinqiC5jkxVWhfjX7vD0Vqv8ACzSGV5DKOx3p3h8QHjtP+Wjz
TPe7UNUQYLwpaPQDxojAgb+R27XBz8ka0MBPxC6nLgb6Kw5nkdzEPsos7T3/1QGdv2hDj5+sSjLZ
v1ppqO0gf8yUnQQLdlv6aG/bD4/hXZU9TyJrpSLmmTRqGIuEa3AJUrm5hZb3mFpqDO4AP+VSPsms
3A4MZnDjWNAR2VyndeJIM8hRer44RyEwlP5As+dfYXxEV2I8aXXvDlLFD+aP4SQoYvOMZNwgsjq6
Bsz3rM2+sbU2LVzg7JcIT29FBUtPSLSfkPAhtZIxlhoCUJVOD5c4kFUNk5v/cFDmNIG2V5kp1Ufd
QUlHBTKRs8+jOouihApbgmfanx///OQh3IKZwolCu06aODa3kl6hCdMKB33gIqo+YM1l1RkO5qOw
aMH/AtNA6XEuHApNeUBtVJ6E5ycaBDguRvlSOg9Bav+iHR/Oi1lWCIpcNPu/pvzkWNjYNolUUmUw
AElGCGAopfhL4p0d6LyNizBAJdok31XzW63L6QSI5qL9E3jElsTjNJw/4RaD2sFTFOdRXUy5d0ZK
ntpPMee7G3gvHtdZMdNSPljolPITrY24or9J64RqpHFD5iNj7WNyMpvo8YwJ3+ZmiTCVCrfYrN13
BQGRwkZfLeb+xY1GSwvyb1cbkXLL6VvJHUENwRiw0WtWt+Wc+H3OF5yiVt6pRpG89znTD20tCkja
YJxdkVS2eAhgbgAp9mUAI+e8ZAmcRAVBWd5qQM5Rgz1R/vUi5J86ZTdV/ZDSa/fiQTdOyC9Y3Nzc
CTsHczgp1Tcvtdy29PyuejLa6uY5rt6DBcRXKZjKR4hoZ+uZ1dgUyHDFEWBnZp38X5hIjXwopIce
AtkziQr4cICThhr+z1sqR7WPqD6uhOGIgGTol8Q38HyO1LOeKb+6MGaHJa7F8mw4NiyHDxK9cUP1
R0x74fALIn8B0oniIcZgpBOpro2yh3EwbrSsDNxoaYryHNzyvJTPv3Jd44zk99zGzRg8wtosV4mx
YNOKIWTfdq2YY6RAYNEry/okjYWxdKjs/fAlzt9TSFBgCsMrDzMy5+zbbN5YDVy9lwxk7Uv8lb9k
poKA423Fj2QI0tkyJlK9j3AGJC5Gf5gkLq4nc84Z1JGU0d0DXhMw+pU2zwROfMcG7EJqDQx6OKvn
heM0QxFSNRSPn+T80JhkOR5eT34TEF/Q3OMAB3GmYuqSeFY1ORyagwxEnx+Qo1fzgeD10ySPQphD
xCMwYDrQNzuGIavG3ENJCQPkaSkgnSIqogurS+SSsM0fxjwY3eRyxWTot6E1F1+GE7f1ciPFYPjQ
jx+33uetn4DPtgiWq5AMjqeiO7n7qDQGFP7ek4O1rbecAcgzA41wgDQhUo7qwORzv2U/z/ECyaeE
0pEBQO92Tg6J+EGel3I5wdYCYh+ZqDrTbGDM4PStmeAYihjlExLt6kZWMTqi9988hhazGxeGI5gS
wfbr4buhsrvw2i++vi+9fkE/Z6i0XYwn9jGCUyie7pJC8OCFbn+OOsNxxaW7sNCS0NvUzJFx/8E6
GvN34DrqwHCFc12vQIf+mzc3nrJ2baRSZO+YLfM024J58uTQL0/xtE+usBQVp+s7ObwUMA162MzI
xqswOa5epgeFhFGdjZQJAJn06zxonl1wpweF0vzIaKXyY773TKQgawCN6qRr8myBH/eP+7S4h8Xe
AsmHXQypouFKIX4YSOg6wGskbURqTEHpXiIJxZ9VG1rQGkcdNa/CnqKUwiOeB6scV6+ACQp7fHXs
kMmdXQvm/VxRcoFSbUn2UrwsN2dU34+1vfG8A3YaQTja/z6N5vTPVxXLii+pt6RA3AiwwkDPrk4B
Sezj6SLQk6foZwFtT8z4oGPR7GPUorbQk8zHQc6l3jHk9R038/mlAR4IrKCtnmZk8jmzcgvNC/tZ
5Z6BKBR1fDZKBvDfRZPokFHecIHY3iie08zJKayDFSyPZNlWhY5OdrWFTgLUM85BykhV94iLySRP
QUqFqt9zFHiAAqwfWHu50FYbFLNPYHj8awTRrs/FB1WRQqLjNHv7PDu42teecJPbUdXaBqcFJbfc
Nc9YBxJSfK7k51OFpwXUAkKJf466G0U/s9jdTjBgmsOkHpqHAz8vVKBdfCzO32A+tFXwfHMeHEH3
khUWcr2SSEO7oIOBuBHQlf+B8gGKLbwsypu04MbkTy4mqNa67h1lPxDOpkCozrBhOG1WLeAneY9e
LGjbk5oWxlZ60SEIdsXqTYjjDUxHybGpgB86dejQZVsooC+IccDwyxKJjro73YldZ5IRtzsVuEEs
vXvLiwXjm6P1NFKUQIZO0UATxOmRNiNjS7vAt3I1pv2M9MCGRDE80A7CGntiDBSSI8Yckqe8p460
+CAyLsmVaV85KOvyb7G08TtHE9VgXl3R1ugmUrQhY0EgTovGEq2ps7v88Y9ujnl0WtculfrbfIw3
25igbGb+ir6SRnzTCg8qwaNaKVkMeFM1BCoaByFLb8aQ4d2KWQN3dpyX6vIGWFTZ0ZeEvwcFpFbg
syPZGGRHF0+SZ0TsCvYKNEX/lfwnZZHt1bECdmM6SBgTg+/iGCrBp4Xy0M57YmBEocFx5widwmU+
2ahLbbrXm/VPlvg4bEpMQKTGyP0UrR4YDL3PbMatL8fUakIZkZRlAhwqWDwyoCr9sKSS0Hj0yqln
NCiRq1uJtTF3U5h6UqMJYz8+omWzELR5+JmDcm3nmEAd+vggR23GwS5GPDX6PHM4dwadY2uhP9SI
2mJifdkmn7H4ESoR0zWgCemNWT70vLNw4T45Ks+NbvX0aJkmxIhNXiAswHbp5Frjd8Yi2hmBeYEs
/caSvvuhnefhpq890Mypr7xdzc4u+IyXPxgbWuuhTf9vRXcXG4OudBW4noz+PUOkJ7mfSQOSoVsk
c4l1mrsliF1yjCObZlGn6OKMQjbg7niWIfhcn7Dwlx0LkJsxrOm0ZtDMiFcPSmF2YQSVa8J0r50W
ncITBmWsiF2XzLuzuvrrxzqB/csTmKuYH98/aOdCrISg5c8Ncd5W/tUHPOKpviL/TEtqMnARpSN0
ywDEYi8Bur+Reze1WUc6fyUnSqC6qeVVZC2I3XtEjamI31Xq5HW+Xyd3+MvElZw9kGP4IoN080On
i0gx34z1Z1pRvs6JaYhlpgzfSqbQkStvM/e/yXQBziGqQ5Xqz1yrUwhJV4rb/CBlVqkUFFRLT6pK
XREyqIMMK3H9jGpuira98/egqrWXHQZiucB1EjwN+s964IEgW9P+j3bg0CsYv/1s+1n9PY/E6J2P
fs5Al85aH+8E1DbbbGdr0/lRL086bKlXGNhXW/M2yiHtUHHGT7ueAC86JI/gPDfoXyW8uE1uHs4o
WJu8DK295E2/FhPLBAP4A0Q1wvh04WfUBgkKY3ZG9scSmrRLOmSybDyFx+GzfP7d9k5/VzXANqqQ
zaJ3hMgNhWVTYFLhXihF44y5mH1NZHbYJksj3Mcz8bAW+JgsOg2NdfUrhawjch+RQVfNGPD4ISH3
ORrsmmw41guJ+VBp4y9hFhnGX98DkoQrJens/lE930wx6sUyIn02n8HSJrvWwuQYtSVRs/mpIZz6
zLIZjhDAR6vBW2DzF2NIlMhrxfPPd2hyrAeUYEAoePq3V6wmprTYQoxZSCU8EA0iPeXdHZZ9VXMN
VrWtMDotGgYySvVGd39k20CNRDaNpXTV/eb77+7gWpzOdEMDhC2v+l4nhNZqqXzVMNqOWPDIai+O
cxLRuJH4/ZxiWGelXWzIjK6ptH1FaFoCt+fdNjDcFZY2KjyCySHrkAhigq1JThnFQsPS1HYB+b7u
wO3uXlVzb+qzYIp+23CcXyBbnOf/O6jAvxN5uwZbRYHnzh+9QoWDkmC1tHDYIEfiQOlY4BrYnIsa
HJQNVdtb7xGAr/YJHyBnl5ZURe7K6uBxXEIy+fQzsWU4oJ4Pg6J5HPvwoGRTUp78BfKgWRoErBuQ
5nk97E0m4SeTpoJcx1xV8PrVgo0hf8cPrbokisK5yUI3h1avN8eF+UZQ3V5OgK6DQZm398un2Gmq
gWQuzpA5gcyP4P0WLTls+Plpy3s9OMzKurb5sHsaKZ983mPhFVbaNxdplsYwZ73tbF2sGj8YcwhX
1TdU2jrTELlbHTlL0fhOFyxT5PopZ0jYLh2O7tJNZZyivJn9HrcjuMOq7MxgnE5wzeNgwcyELif8
ayAejzg9lii+cTVGQzgVnbdm+YzOXKy28J4/UntmrKZJvgEnP2zpE7LfDqABGRwYYSdyQEwcI1uR
tmZXHffPIEFml93nFlRzn9zMGpQGqNh6cwa5StHKPbpArbIDAmb8WMvD+0QATb/2239Q1K4wpzIK
Kdp6UnOY2H/IyLiNKKPYJL7V2y/qp6m35nx4mP/QPdxKywwjhldcrlMVKay1dF+gZdVpx53sxcIo
aWGlF6jK3xgOShGmh6pw5ezrjTX1Kmob+UmWyDvyL1eaxLAC5+VYKnqBWuq2zg5fU1Flsx4EQQCG
S6mjVDBFtVZDCQtQf6yuDNlFwolHVgaMWuwuItD5ndClRY+z31Om5Ts2NKHN+lfjZVTt/917Y3Oz
ngoPZps7cEH4a2aSliZnJI004kqY1/E/zyYywxjjBhCyZrsu8rI/OeX5Gw7iBOq8+2tdh9de4ESG
Yjta+pxmI0fOrvPUxmHh2IyFJ8vsM9eB9wiPbKJcijso7Bv5znxlAQUgRT09BfElJVc8TP8qRs7q
uk8Jd2OIGG6kpB3ZN5uSicbY1A0ojnu3HcXXRwXnTVhpj6ILnHhU0qVTQMutOXGndmDiAZ1GQfYF
Rt/L/YrX3ZUSOdDKK1OrdxyMtEr8P5gS58PY+oqKLiDDgbWOyNnrxa75QVTzCY6lYwQBa1pH2Xja
zAVwp5i50IEv1vEx67o8dd3gOcgzS344hb8frh02MFGPoLOL/EgUgmp9OFPrI+K2IEeuZM1JV/+U
Q4T+s7CoVG7K9XNrIagA4hgeVEW4A14gP67Vpkr8c5hcQ6QMMghgNKekHNBS6nR6Xb7SKYSUOEjS
XaFKcdjeGxEukdBFBJAn+2YF+H50hIJdOnGotYXE8VBhC28H+zfAdU3XNYHbuLZ13QU5/amNFnOG
YQsKvMzNUMr1IxLvY5lIr3jVMJWyBg13KXK+kVR1UDiKasZvOPWLj0HElxwTKfkSIabNVq0MDUKx
/EcAp/6BNX4gPDl/OzJJbt6f92/2DuDhK+b7+OaeldzshxF6kWmwholT0KQ1YT5dyrTuVmgvWu1K
Z6hxkxcsKnV6SujH0J3Ff9aoWHjKzsrat0mSsTA1YtlP6+DH6P8GBipBIBMEKVSDpBStbfQCxD88
Nd94ZVK5aqmkZD+x28hp4B9nBc/EA56QvfmgBB5Pac5RThcjkkFHakO40sHPH5PMpGCHuE6qrYtZ
A1BHYRC6G4fZnd8+notMLIgMmgM0RSye3iG7+nyDM10xnZcuQ7w6MEh62ywDCCBNDuqFHtwNXwK3
WdPg/cLS2eWAWQgrb3cWO8zrBNlFsDKF8l9S74yRKsSLAX5fZJp6A21Bly/gYH/je6Rcqb15ahXn
FKSVx5ep26G+eoT+gAE9JSUZFH/qDNai0K1OF93cICrGSrDTg07xUQGSKOaPOqP1SwxYZVC9gGEr
xEu2A8nPVcptJI60xzXDa+NKaHNRt9YpP0e/BSPJ2DFPLqy4+cEEzvxGE3aDLNFxIk4ac2aqdaID
iqsYX1xdHbUVC1cDOXl2MuZPfJ5q5Of6BZxyu69znhlivBj6AXGswYi8TYk3U5mP/Qkdz71QsGPQ
aLuSaIlTPivg7aRVRs6nW8U02gplpeN0urxf0TYoQrZ5gBsVOK+wMbEcgY+XkKjovsQWP5L5M0Nw
RTb6MPFnNIEuEoy/zAUm48tdErNJRtN7adaWG0lSK8CeSrDaUyJt7hZ/nuZDeYkUxDGOuySXmV2d
EQ9axN54E6thCe8c7+tG1ywbAbYiX2Ka5lljm918XjGD69Z1ZHZ6IPKDcMvzWSTBxPXS9OBWJurv
HQc4UKlKj6q5AZgmJ3vaiADZZO7+8aal27jK2LTRGmjdIdnOIeZx1P2j4g7pM/k8f/2gbh6/YtAf
LKqg2lrISvbQ2yw9Oe4kp4tzmWTeJzZ2RzWPPaMv2DwrCp2yRcKqRT0dIVHoDURIALOyb0HLXLZx
m6OPwLv4kadKnVrv+L5zO9PPjMoNU6CzKPm1NwkfP9dj1wVXfSQyKc9HEqU9y5HkDUWqMg7PmXHP
bCzfyZKLEtNcAz8XSY2SqhDOVR2UFGjC2QKCPZafZXfTFC7OfWlOwDkEzOZLVSjE6d1+X7EBj2Sr
kIc0zSqrXO2thK2JWnAF5YVww1JTo3Hy8TuApeXPGysSomoOU2gPxYpngMqlU598IV0dMtn/POZr
R0vyVK5LMRTyZFgqefz4FBu1Lf4dhbiSTt4TjZZgR1WoPETQtP7Osjaa0lrLu2cumyB1MLZ/5cfn
w5c9mEpHRiAayR7I732qBApEmwGRJH0Ur/uZFQH12wFrxv5fmqLm/eqT9W+DxvZMrQE/l6QNdarB
Pz9RytwsXTMbi6rZKAd4CF57y49lLsgGx6FiGmTWI+R38iiTrta6eFxiIE7BMjPjSsXXtyHWp6Mi
MW18aP1bkZtNFBUt0SgKQBsjdcpiw8v/pxGJUyQoyW71c7buiJHbvgdlpistC/15adU7Yd/AO+Ld
Qby2rUm2jDx9erwDXC10dxHl+PG1sg1VZarZy0Z5Nv0eMYRObfZ6FmXGAR0Mlt9dz9t54NVewfJS
7BbR1mZHuDWf95FdiQAfDDh3CrmJE/C5pQcxjTyYAYcaH/ks27dFOyx6LVxL0zE2cjDy31mxzs+y
0GSFBWC/s3j29Ydpcqna4p6evwK7zC2Eg9faIFpupZdeg/NQoyR7agyM2S5NpDAhrFL1GStTN9w4
T1xCRroWWDkzXG78L/EHbGry/qdDCeZJPofPR6P5zDb8N9PZa4J6oH3IbmL0AZqqa+G4cQfq8QVn
ypAV0xP3C53omG/CEUOBotbfIeB9vbC7QNMUaEUdaSoc1ziFM+NrTX5EY5Yg93qnnc1Qr3zbNZr3
yFWMX2MIyRuKr2BIu3OZ/IzuHNMCH/jsg3Dj6aL0rU0E1eqNL+mCTHi4HZbEyZfZK7UCU6KBUc9k
MWEHO738IXAijFkR73cq051X/ZhWkN8kmT0v3JatxChq3StTRjbIlVK0rxRijL/tBdc/aL0xS5XL
qwdeZKcZJ1EQqEjYo0XfacCtS3pPsrAyhFZ4yEmO9qjQrcK7liwIfunQ7/5QtVVVKpm7Ww3toIsp
VVqkRxZJni+nD+7T+VH/8icetAzqsDUKUCozKi2svOzA50FHT9oEGFL3KPe4/owgh2qyLIT945P1
FqVkIaeVGtJTlmpieXWltb+KhJbP1c9qZ8HYqxxPR/xGAMeRkAY3BW9bplP1Od1PoGzZKSBPldQr
9AA9PC5DiNoNYykXYc/ACuhuZ2J4O14rZrHP3us2ZBA3eNMD2ZT90MOo+4STk1oGaDA48guB6Ys1
9Il3jQyvan54whBOQFil27Q7F4eeJeAEk5c7cVt8sdtUhaBLTUXVrEqWYu0pTjWRS+iisp5kuGUF
dkb+elv7WfUOMp5rGPKdZUKDcrTYsv9FQyNET63S/gfqmnZIH0AuynjBS5fKcyUEf7P6mOoOHBKi
9kHIvp/y7uv0IbOQC3YK2WF6UIyZzr5sKZHd6I02qoZIaR+EEmUoJwAPaP1F1sRA2Sac4up42LB2
T+Gshqq5tz9K+8+Kxowx3ykjaPjNRGZuXtTRN6I3UPH71Sw5OfCFvY92a6JnVXLQX9fzdEjUb6MP
eK4tftb0iX1vnCrdDIrhKpbhaVYIJ6lIDq1/YEym8yxEG/nb/1D5HR781jtTlODom0w4r+FIY8de
m56z0XP8j43Qy2pvVXRAk5wE+13gsuD/zst/dPFt522ntBKzrY8NL9tjY2GQGL4Ful/t2xhJ8HKK
3/i6PCZCLKxgmByDw6nXK+qWFtGWjc3QEVm4gF0nfegK3o9Qm2ATWCU3QV3v3jE4VImZ7+3e1jp3
Sa0oUa+Hj1Qq5rMhemLL4Ugvo7Wk3G8Vw5sdjut4iUvLWIgROKcnX8wENk+xQLrv6abVpu/p7wdm
EJ/G8CE4rhlyJ8xdyI5xgNHfsAZEmvxxD6SqOpMhS89W7ZJRILrx9bgsHyJW/t8CvhzdQki6I2Z2
qMtsjC6HCcPNaXvmxs3EOGRwYJ5e101IpkbuSjfQ3tjOoxfc5R+Zeskn6qzElarhJRP4jnYHH87n
tO3kp/2VXXz6PkmqATtS062iUNMuiOnY/FluIAMHGnTogxk1juuRjJNcqsEWcNfpNpOW9GeZXcPH
i5iSI4vKEDqaB8tE/poualc47Uu+JuhttObviOb7QF90LFFfgmHKTr83S9nLA+QUinDUN3yqcnr0
Fp6rTxMHyUCmPcpqqwXvINPFzIHDbeuRQSNOJW0tz5DVNo9CcgYeJn5Gsk763+D4XMTLnAVaAQmD
r4Y0UXPq6jJeFgVyePGYxP2ylY0otheMmZetkSnQX/WN05lOxyIPPFUlSnwyYkmu1NVqc3CQVuwQ
j86qihigDeGCf5yy4+p6wJInZL6hYtDCr0VgDkRnro+jy6FMLT+HTm/uLRhE9mIQ+9ZMOsTCbtv2
ikLyhnD40d3to1s3mugJJ2wJ79lyXFNFfJj0u//+Cij14GP2CCMfKIrF6OLumh/n+bhQqZz/rJOS
mkJpi0o2Xd2ph2/D9nlwuGkcjfRjABq1D732HN2E77oSIS1WrYfw4Lbh1kB7/2Tq1bePZsYpD3Mn
IHyjEJulJB+v/VlWuT5s95bFXlX+NED2CdwLP+d76Zps1Y2RtoAdz5iXGdvIwUw4yHeUmWtUmUBg
kE1s209yDujsaw2hQzO7Kj96l71mOcK8VVjekepJH24JBg+DxSIGTr88IgRxGTaZT4hYGataWk/i
n6N6iPy+cXRlQlTloKIWm5dQnIc2CeKo7bgrHj4S1RWIQYWzO5nB4XUqnKskkxTSzL9TJnGS3spJ
HKUdN6HRkNUR7/Z05ucYrIKG93XsT1BJn7Ld9JEzf3PgiUCgh7fO+h30+yyc0Y+ebcoHVZWyvnDM
qCnXjrXMAhKUW7+tGE/N8j6nZoTkmQ3zZ2EpwgjC0YbJHNVjINoryggMoc1HfNBejJBaU7qdXJQq
8ikIZdIVHOIwcXZX2Wd2tkH39FfksLtsEDO2deQKs9dHLtt6nggc5kHYtxBXwPbzNjuq+JWXN7x2
9JVNFwBQEurzbgkpdT0dSO3HgiiCw9d+qQ8CCjFY2VEYjbttUApetxMLcGT1trP1Pb0l4wTJt8kX
anb+XHcIKjZFuw1zJBXCIygq1/16GaMeb0sA9W0Ry5E+UaIZkbtxDMC+S9whPt80RDVWG6RKcghv
vHXe5pkfrczA4bl8r9mOKzawwIGrA8SU9BLnW3rzmgRaaL047jyduvZZXbtvtBmxE4HAkgTQWRnQ
C7O137GDucZIvQZG/m2149o6hO4WmBQfG15otEduIAhflAFbA9OnXWa+YH63iwaS/DHeMWKoZ9lv
shijweL3ve3iguPoXMD3wtauraddjyPRjKQgJ4Y2AVdWMkZXpTTV1fGTaInlxyYoOiAoduXNGvRd
8BqTTS/Sz0u3sgoTdH+HCf1BZvileFkAzJFtJlrcenMQ2Zzj0OWAPv2ssjHFW92ecSZbZYUFriBp
TahqRizmWovrSE5ab9yQQytTKsUq0XmGw4Twg306UN5OEYNKkJ5wz5U3CxjYj6Uw24rHghsTIo4l
f8n3UnIDGzFADPuGs7xYZBhde2/ZndOnohpQSGF7pJMvqINwBsXMy/L/uUG6gCz8JrLABMZGs1Lb
+fuwPqFW7q5dqQxlcWO5oylZ/QWXV8q5OFBKtudgdIFEpLbbtpxg7/nqvCaNVerHuwcJ9a7I+se7
BOi7eGKleyRrQnpv4B8UQcaJamH4Y9/eZmsQKGV1UUMbeoRFlzEmztJCBlORBrSGy4RCcHEvuFQ+
OrF9EGZvVeqGDqaysXNmRfMisPjBGQyA5zJm8MxQw7jrcVIRtotImtpPAd9xeKOJlZCH+kMvkYUw
I1xhufZJerWE8ePRmKbDUI5dxAz/wtUps4NpoWNJdO597d7V4xH9V4a5/9q7/tVFyIbpr85pCGmq
5o5+XbE7dsMCN+wAwN3H7VaR/dYWIH32If8TuSmzcWDyju/ml/dgvM7HZTg1OtjV2JG79ro0NRYR
9Is3RHrbVVi1OsLg+lpeQYzFyVyZm/2sHwKA4hEKSRt0EDv007q/3PRN6A8+e4mK1KKowabRcYIh
iX5GqQCQMcDxbT5A4hVj2L0TeUSl4eD1Fvh/HYErMr0I8vB+pwm7wt/nGFvDw2D+Snew7EBc1ARj
KMjqNfTpsTQNndt/Njz+/gpeMgdM6fupDDzxj92EzJiAn6z6MRHG6fstCddBnDOTupJjwr0xcFt6
QEzmva8V4VIxD/xFlwoiHC1/nce8YPQo+IwjpLNFDIcGQIF1Aj2prOYpGcRs9R9laWwMgceFWUV4
xXyht85eV94kX/qjKWeYjTf84IyLjbcufXeLl8MSkH6R4M+PpwP7yxNThUEyywNvNM4/9nQdXOWQ
PGUxL1H+tfv4qoeObY5NlnjeYtPa9S6kMHMSfS7S11opoDUchTWEdeEOsr8/TMhQ3alanrOyJ7vQ
43A+yWH9Ubrv4sB0Z5KE2fopmIQED1uOB3L04FBQ14DiQqdAXruatcK0J3JoTv2fzBJ5zfvGWoZe
FM/vA17hp8a3+WtczcjN/mPCHCbrjixjEcoRBYKieouMhWYeB2NtzKVt37Sit8Gjyxmfqym0hwZv
Ze3nu2iu0C1qUMTH9CKhFwnXdHlHD8PUT2N6b1j5+r0oq0wIp5cr0kyNfkggeTQhJHX77989xmMw
YNh+el+O6xU8yTJMpUZDhj7Y21mDI1zyst3XEqIfHlnUNm4qpqpTOQO7uUPjNW9839if3+kYhBY9
adAvomYqT/MesYGn3FDyeZCpk6zaYZfWKrorhmK7GvH5LGFvBaPKusUfeR5YJYntYSqq2sSjYMQW
OgyJ12MKdKP36Q0n6iQUmI2NFmfkTaZnJc7zvOJNNCMD+/MKOMhl6JsfH1g++OStLkUvArFA5AQM
NkaJo2UjigdXgVrfoZVhb6ghxwkxIUZn6wbPOqpDLZ2Tkqg/vcwK/loYl0aLy4GGL/O7InNmPG8q
ZbISSMiWSIprB+ReBltyCpDHYrETXtTvyzaSjkYLpNC2lhLXhCc7pUL3hJbx2tWf0uF6oj+/M15L
hC4DbhD1LRHJvrEaZi1Kwdr6KpaZYraHDt7nEg1Q5wbVx6GJhuI2RkdvxvS4AAukRf6eKL8twCC1
IbZetTvLpV5+NS+Au4haCeDQEIIgJGonNAyI5h/ax+okJuyIJEAWB9zD3keLY5BTKCKy+FTo8ZQf
HMVXgcnB79v/kuCa7kAaYMj+Sf/lPXK8YUIweQYpgFJLbNcxG/GvJpDJnn3BjKcidaEBeWbo8t8F
LxKbwVXoHe51C7Fsl9AFgEcXinf3EdLqslsLCSH2qC7hblkHAhRcIz+cNNON8Hwx1++ovWXqujz1
Bsu54THdafHpQN3C3Qbeklj93vLA2wT4pPpU9ZtY7JxBG/ozAatRnykHzeizqpDrq4FC2o44W4U6
0lsZLShyj3hNLKXinR2d2H4DybrJzfnj9EffjCjZjL5xdBxTuCsS3SrgD8TeNDfl40T9If5991MS
UjtqGOnDBatYKqFJZ4QkdVnCicF6hQjgGHSCZAOKAwp25SzV+RfE9y+L/33DgDS2OnZxB0o9zPxl
3L+yaYhXJNqJy/tD3+X3kHqwPuSAIa3AhF8GpBAD4nbtjZyaT2kKOMKfE06IZWECL6lzaYS/BU2K
yTR9GO3Xx1KwZfeafpa1A6S6vZyBMTcXtAt2BlcbRuTsNgFaKYiDS487UFsxGk9W+2wksqcFV++h
9vldyrmAPogy9HTeN2KCB1yjbFeRQ1RlK9vWZY+t6B7HbzCPsDaUChvccwFlKyrc51VLowX3JEJJ
Zba7Ur5yIo3YnaR/j+4vvHlAGeN2F/M5mKMjjyQrZoPSjXDQqt6dAKzL6/X5EpoYgJoEHvSEPIDX
eMtk0g+Hgiks1Mum4R/F8HOJW8mJHzwhrVgGehNtMo4HkAtQs/Gaog6cFJWIXPu9a20EcJV14V/p
esZx6lFVWWY55OBtThg56na8GNOAabkLN/QYbPAnJPY+WYffENnX+l8yhHXWb1FsX479oUDfY0On
OWH52Hzmahm/PwHlNDtRr7yMQ1xVxYyUcedmAYR4NP02cyFdF682PsLSrZyV77vW6gGfUFz4VbWv
S+fb8coeVC46V8F32BnSg42M/N4HSRl0M8GxNxYEIs0QsJw6lMt6IBg7GX1IMhfq2I3xMj72MzmC
780O2eLjoHc6Bnp0XGdtLTCi2qGxhhsB88MMUkFwhHHzyZwPldVdw5eMK0ZT2My/wmtEbhttA4Lm
1Nwhp8ezOCbSAMYP0PcMcS//KdaLztPEXAmIzhYZeyroGY3PafZ/egrUJLVRurylw0gc7sROCi8N
+G1/6SiUFqEYktDEqNP2bAfxWa4RaZCUryO72l48h/DQ7ajNIwUJMPTlYM2eDIiLRXpFPu2TZur/
BYYWTx4t6t6t6Gsdid90qype6XaCeW/0TVzeyq2w1nqrr++30jWPI7XcuhYTrkB6r98GpXwVC6Tb
WlQGqZQCFw3qvwh9VYflg0DNwxSpGDsaB5DubyHnoJ0q2NQNLC3lbZ3ve696Ea9G1NzyyZc/uPzT
58w+WdYQ/5l8U4tcybZJsjAQWIB5OwwGp7HmchjzFzIv6yz9Jg3083i62jL1AR/ZpR9fUuBCuPzn
D/186bmtktkFOAdTCw4Vr1gST1KGo2rUFV3dQ0dPyb87q1U73V5xWbjUVywNIU6shsiH4o1A0eni
emyJdAy4l5gPJUzcp04NzURP8cBT6+9yCrQeyCheDYfu/LZtz9PfBYDIJ3Oh9OOyhInd7llBffL9
JgvXaJN4Ea1Jr8qj99ULnIe1Z8DzJ6rcuv0DtSDAJmPqEKkmBYHv8M9of6krAUneLp47u2KTJgem
hB4Ec435rGLxaGxnh2TQqkz1VHoPpWdAkudCpepYX9WTyEXxWh+8hoklW+X4mjinJuwDfIM8Nx77
VzocbVuL2bIAIFMW5sSTlZdiKfzlh1OUuZn1YSozfSuP6tj3ZufcYyhD1iwfGZg2tv1x+KoTzenU
0NIGkQ7zKpPTBFPKV/K0tisoKdMsBLffBD7f+iuN2dB7zjmHGhSGN5XPuJtEWjXzK149GMBlWmI6
vM/+e8ilavQMx2zbXWlfgTFBwg+lIqqTCxwLhRDroLI7zn0G6y1JCEKOV1JiiUc1Cshj/dB0D5Z7
bt9E2ZZgoBFOYxaiH/V4PcrQ6WAo3kynJkGecvOJnlpKyaBTGadTrx6ZF7LS6edbutz1KD3ZvRIh
pSfKnc+vLiV/IsV+rROeO41qts2r6q0LR27PZei9bbwPJ2mnXTwPNoqA2rMSDtjd+jTU26LQfSKz
hRRcnMS/jSCYAGeanr1ULNiVaYRYCbveZkQqjm/x7+XGByQFgVSt+Z7PpceUJ6HOaSwn5qu4WJs3
Y5iv25pW+OIlqPpvnOoPgV3Km9sLEKFpd+5ILmmz9SP5fI+LM0JCLpzT+vMv2IjndNvZOPd+bg+r
OKSDQjp9HPoolZgbGIo5C8NJXhqhgAeCqrMCLyEmqefFT8OFy+UNFN2weLnt/dMyXtmjsyyh09wA
IoDi4In7iCdw0yu7GXD8/QvRcc+MMTSx2DQBC40IpDROcmF8VUnCogfN7iaFuYEvnMCqcw1NO2vf
YDUPB1JST+rI8vaeIp32+ejBATPMvZrQ/hz5kkCJOW7NTy7mRYZRk9hv5vQr9QVZj67OMJpjduRa
bACjwimUGyjWrKkFf4KMNIP/czaQWBbww6xrLcS2KtgR7MfCzwBJ6zJloeJ8j0XEiNqoXZt/B+cL
eaES/B0a+pfoAQJJ6zuxL+t7wwppM2PXm5sEu4HgnLJAMaWqo0puMZHX7CbUJilhhIN7bWDQ1ss9
4hFCNEHoMPHXIewDntPfo4eo932RSdnBy9UKNUovNagJtltp1a4MhbP9ezU4Ue7WIe9AlCsmlAEt
tQJAk1KldkKjit5fOqBeFkYEj2xA0BcU6vtZ5ceUuDYE0taB8QwaptIMPXindoMdDtvTlXu5C0IZ
ZccvdVMBaE5QJPzKMJWp2QVlYK49ly0vbVOiEseyoUjJK3LuqHNrObc4JrKhhDaGe9OImf7aDd9X
wPvnlCa43zCQkAw6aDs2CQKH6sM00rwxbLe19dv3ik5LnmGOPz0VhFVwPS4feo5jhIaokbujh8pp
gSU8oo9XGAXwQUI5qNMvKK8Cn6LHArxx+2d4Yg+ZjJdvUOiwdOE+ZOFvy6rMdcOcwLhXfGMIhR4G
OkBzgWOTmprMHmO88mAm2miiirsJIg6d/D78jbgrdVNatBV+Nz1gVJvhFZ64OmDT80YU6WJnX55V
CyKHL6oqS2S/uH186hjG5s1lVaAxYdWdhQbe8d0vbvcBpXhwASa0YYbuIrLb5evtBKra07BEzfsb
Tn/L0pHRBl0wdRimqwsJRUUf1e6f/AfnfCj0OOu+F0xm0Rik06lfGTU7w7gnqFQ51OHu+/xD4vE6
sgxttclA9SU75KclNZsXLGGcqDEE4ypvEK6OGaDCCT9v/6l7Xdil6gxqGDjjQI6DRBzWciBcM9kt
G+3Wu+1vdZG5EeiSit7cyPzsN5/JoyRh9K3mEdy4PAAT7yg1q5c3KpQFrz6RQaXY6BK0ptIhmthH
5ncJszfxNa2u5O97C8V90GCC+nKYDBjbHjTvUN4Omabzu9EpAms20ZigH6b+AAGG8Cw0qhViFmcE
ewd/+Pu3xiYtZdmWF8c6thUIA6VHq+cQBIWDyO5IEgxv/Z5hEDG70XvwYEj+4KRZCkREcg41mJiH
jcitLvBffvIXKcHL7ZhRyagepPxVe61yGcwKkWAGxBJloe/jlBojQwnR8dU4Hc8tGkWNHVX4WJ/R
+LuslKcNNbsnfaGbhPXv3MsQm3f4Vb1JnEF5MfpGA4eR92Z5U3M/xkNPM1946ObXTSon/JhUEeRm
QaUM76Bf024EAxU5j5rPXjqRUfTkIgcVSg/1+5XkjY1vYV0wbZxAL60nPKUQLU6HOWw66H708Myf
tdUqwKiciuGsz3JaptIcEeF2VRzDvedZ+jEcbbMZmdgX34jKTok/8G3RFlaI9yxxG8WyWLpEuovj
oKkOVZ5nXEqi++ifs/2eztkkF8fLW9ogg04q90U/Fa9iw7bEP1B5r+8XTyG/lMRLHd71GxI1/S9S
Y4IFH7ATPqUq0+e9dSUx6Q/Bop9fQL+lLIZhbtX1+oCHBoy9yzovXrc7nrZZoK6g8H2zUpOgiXfx
PND9hzCPB3nRDjdyXmWB7bt3JSXy3s6tZf2wQRYfUYxXiINN1DlLvKUbE27r8WTEF5htDj5HOz+D
1sZzoztqXBJLRHR62G5zJPsqQN6YQGlaJ6d3JIenkZ01R/A4igra+iHfzPhyzY29OaAIp1MB6KZf
sztJRRpi7vPk0FGPp76mr7TKt1uwfjmjITEZ2pNChZYDMvCRzdqXU9VuWG8EkjXGtOWK4rmHavGa
iIzbx9r5triCh3gfV4K5WmZBdhEvKr4YgzT841hBOO5RfFyVPmmPpWwFeAun+UaSthB4xqH4VkTv
tmJ7ujfEbT5baqzoBu2pMcQbT6VGuInP5p8Mx29M8ytL1BfimCuv58SkdbcHlfAOVYyvGvzWEcPV
Bc9fWxJZ3kAbcA3xOKoM4hqOe+msXRnm1dwl2tHcpB1aYVvHWzOLMKfXqF9wDKCGRjVfJ3kNPFDw
uz78WEUeqQOgLZJmUEyxAYsqat0A5AtO/I77fci2fvWrKyWHDnVb3k9DqU6Kq5CSRpyvu0QYyji/
yPW9ebcnb68Iompu0+kQsG5+7fLLVR798Kb0IkKN9JBghCz+z1eOp8hAkU2NCTWymYqHi9eqFTjy
kfqJBpkYeTYLo7fMU0f9iVPm8PWyQPXWC0f7lr0+aTrCQEQxvCjDxle0UTnZdZSC2uiA09wQKu+5
a4RhIfMHrn//9WxMmYdAMz3boub6x6uL9WirNrXCvHCk+wK5BlxwxqOZ2ujSVdDNGh2UXw/h/qpk
zJ6RwvJxm8ZcTNHHz/9P6raHvPTww3ZNXXIRLVUpzuXful6jiGtoCK5yJ5+UoIFUFEavf4/g0vhX
u95lMP21znLdrAbFUtKbVXo8TfjFfJJZfcWO0wQniqwKKuFEx1kk9qjtV9katWjCQtFSJJRBTt9w
WE1/x/rlvtG6ud4cWkBuTOuaoy9gJdWxD8zD8xVjZnq3i5nyLknER4Eq43VZJdvm2jhpnto+3cP/
hB+27BfEqTms6rS8xhjcBSWbbtOnLJbLeCRCeVIWOpoCYfHKlkbCeqXH81+Ezxch14NH/d06CQTW
wBDTp42IqogtrWN7oIglL2+SifC+omGubySS+IIGeN4HxwRsZ77G4A446JZa3DHV5ZDJY9DRkxbX
1lg6vm1AjO7A7CGHXM3n2wkfUVTH3cPW+dMieLzpI0MbSebmFvptmHml9EQpMCTygy4usQaK9doq
0YTbKQa1aEXTUtHsRs4cdiC0KEZ9Rmw0qGhiq7Oo0W10FySNKjskjmPrrLXAM4JyfoRlijUUjCp4
A9qMr32/hV+hCkx5ThU+H3wjfHICh/oiSolmccA0Od0bq151Sl6LdcdfAWfN4fwzi8SGr9E0mkf1
dgs1J4JpSZZzHQw9jYemAtUjpoGadq4o7IoLvh3jdVu2AjJf+XGU53o/WoPiCOcgSodo+KOOB4gk
0pLZVw0ZoCY3z7kiNN2/ACXvbPF/Xbr1XVFeQSp2vksCxJQDRN2QrwU83NoO+shN7zp+XLBWvPm8
aMmQgNT0YnVusc2dXQRy20SPXtxuJ+frfh5YVKV3/GztlwCF2wOQXal5q7jHNC7NjjFn0wBNF832
U9peQgIawAu2deZSAGaImO54+KfoTYyXDjSLiUpZyi5mbRZXGdm777niO2JZgtUU5FKIjFfQCIXA
KDsD0lTVXcCSbfL9WfjuAe46mxoUa9lCigajIbKU9g/tlEPAR6NK3va7sl66DX8Iu5BoDuYo5wdw
KYlHhDlm1pI7Z9BlkH9EbUwK9woa+YuaUzIduOmy1iOdM9gyC3KJlNbMeSKskY04w2aYeeZk1ioB
ovuJm0KkTlfzKPCT51sE6aDCa3GPSysytu66+0aB4nznQgstnGTrIlbLoSd0ghfLSxkg91+Snocb
TZqh7k3+sJGutevJm0qIBQ7ib4G4x1FY9V9PUyQMAy4uItn1L+Cq8Cc8ybzDa77FhQL9OUDuMEjS
mPNAtXuH2XSTKBjjj7vFiNjbIOB40zkiUnYYSldURdoTxXfq4wrAVnEkTyJlPtRjcDuHe+aV/Mfo
rZfxLEfAocObmyZ0WU52t08yFmupR7r5G3ITXGP+qHyrqbqeKOrhjLF665R4n7DR+BHLUr5S7fNv
+1+ehJat4FI1+1lxYI6QlcS2Y4qcLD7qRaJ3hp8kaDSS17Vd3X/yvo/PfbpjsIVtxBqKdhjIXhma
JqwwI63oU5BxNCzOa/6TG3Pd3ZvI92YPFaecigEu1zRAjzslJWJuCzVmbpQCDQbGI/mIaw8DpLL3
5Z2Yt3I759YbwbZdxIZ0LJgRQaM5wvCXXDe7KcDCtvhZWn07MyvG0FXiQnNJbwyZDxD5xJcrMxP0
iD0zqTS51kh0T9s7l+dbV6A+GQ9VE2wnrGPUrbtFFqKcVqLqx/9rOCpnNQdGRDieTdt7iU9HsyNG
x8MP9gtFTwAYF6TqMIcpu7h3eE2irewMVN71cZTWL67+oFzmbryrlI6eT9DNN6w8qR67m3/LujZ6
xrMC4WQTJlfOaRaSOH+QqE7jpnB5mbApCqK+Kg5+R/32//BzMVWJlSvqrCp+5PORkmTEhHNgL8+x
ELyvdBzSrHGm3P41xhgSza3Sy4olTNpDYMR/FrSsIIR13RoVs4G8wDvZ7Gr7DxO+qjCVq9+/Pl9b
RZI2o+fWJfPQybE0ZENVSlD++L7lSlaD8o8ToC+RLIj1zm69Vdhu9qwZRZ4FTkx9F4qVWkWIxEoq
Gt0Zzn5JJ56BUT92DafrnkQEPCJO/J9KFBdOtkp8RCE7A+zu04kZpAxY0Es7N//9q5nwCjLaydhq
cH4APzRHkh95KW7jQTpTmxdplX6gwtKObZmXwbcb3s8/RnXlnLcU62shVe4E+DskENQKgfVeL7n8
J263sA3vIECy24C4j37tEUlSCvHkMjMtXthy9FC7YdHj/afEv89cw4/0DIOUl94UZuTEB/P8MrCf
L7CF+Ul5Is2hfB+WuhcJgxEThQJ4MU5Qd2nzV1nR7pD+wjDyS0ZN/yhl2tMRFpQmZ/g+lwM9a8YH
I5adrfhMynjFjN6Gz7H6gu5kgulRAQW5/1N7VpqquSRcOqhXz/6w1/EJtyisrest3ysLISy+doNZ
pStif/HO8+fs16xxGrgMTnvuUCyB4+JgopIQfAUDkuyCm/IAM7taOZXanZATH6EskRrGtp4Oja2L
pM3ezEn53H/ikQ6229gk7i393bVb28v7g1kbNxWIIzjFroXUv2Vi6p3qaei6XGVPKufqpH4g2va9
g6/8I1xRzvYF/e2G5WU3/y1+ym2B6PXd4AC3rYi0Ox06bzfPam9OnA73Yr0BvCoge9qdHORoREnI
+SSNRN4MPHaHzKOhpWbrOb5zN3hh90896O7vl9rTobwylbPZjNDzaUG5R1AhTxOOu9JsU1uk2JPZ
pJFyrisxVdlOVjFLc1mBCEVnkeeJT96G3zjA9J+5x5C1Xt1vqmniBaspsp7V4IdsFA6hMmnilLFJ
6jx3AXEhHJy7TFOvIvLw2t3btKcucFo+/x3ysX9yB8sJZH4+nUNsGAZBvqNPMWUE6JH608d6JhG8
2z/IdzpVokElM0IHxtKLgd6s4YNuMkgqlAU8pXt7kX889Ra1bFBkYMc/tm7jKFZYl4dlSgcPUCfm
xZ8D0F/d0kr3c4pXRVdjudrjibD2lYF48hHH1FGK5Xud2PRUqDSt2uuXFOSKwU/6G8Un/S6ifIGX
9VFIFG6byZrMkjq7GLIwlrqXqivqb3Osy1GRb59OYiS9SWI8dy7A8aaWy7VHqLF7KGG1GjBR/Vj4
g6M6P4hM47s+HNWSa9LA2zjxGHSLdnX2QKT6JBdiSK/dUD/MJgipaBXoXJjETwLQ6pgMVOrKdDxv
WJ4LKvXKrLWvixTjuQCKrgK3hwtby59Aw2+cI91xW5sa31qhyU58v1/DW/IbDDrObEcQFNXpMnsf
D92WyAEhp9J30OFdIRa8umVkyB4JMPhh1O4tWFM1Z7Z0cjsAC2iKmQDyWlQrd82Czvy3ZSggwwET
mxr3S4DSrgpUJgsurtjPOV4o9KQDeDRvpbzfnkY5IDuuVMcRNYRdmYVP+9IWGW7Gjq49RT20mcGD
VY01+kl2nvxLJg5xRhol3pEwyzZ6rsCmV4oC0yz4vjWiahGT5AiVaX8OwclFnofa5KNswDrawWV7
M2TD+xV8FiZUsw7rUVzvlNxNHpukgJNIRDGSDrEHYw5kCDAazoAz1dFQ0ZvzKEvLQEWzSLQYPywA
73c9himVgOjbTie2v3VJclZ+sicOULdhYdVkxAYXdQMMBuELtcVdzG31TUpjjGkELvft09WP0Fgb
nQf5CwFS+kqF8MII1KVIZn9okCEl7USehZ/i3z2nmGSnzx6bl0KIw7zlmuj7N3T0YLyDuE+rXWT9
x2IYlxzuWrHtX17gr4HldarU2sfStBo6esl27+Zd73BTLq75Ix0fWwWTh83/pWg7UkZF+bXu//Q2
xpeH45EGO6cZTXm2u7j46r7W3X95gnE4j3F+2vrxk82Vo/wjDN455bkoO89ttOdTbV5QRqRotEyd
dJIt5XubbD5/vIno9XmvcBCQtJ1oJ4IsnRYsn2+IWOPaQkWSKgo5/YYe2DbNEAWY5pB1jmerNR8B
H2UwZnKecfXJcZulDUK8SSrQlE7R5PvJkZTW/+4ocz6VU0uC/Hd8USB2Xf8nQgadwDQy7isg/H5w
txpZHMknia02uJN7wQpCc5DUMoT7OvmHuxpuiHhIgeXzrxIohCv6+WueQz2eEa78oq7UM0sLIIrG
N6rRpEcQVfiQr02q9ckyioQAx4bsHn8KxUu/glCAIevlwDkCjYQ7jVHj1ljyAnZ1jJJxoZFDKzcd
20PoVz2dPCNen+LqitoJeQPMfodYaSeL2LsLcecMbhBdrJ4x26iJB22DVQ5+n6zsgzIrExHWhEF3
89wBIFEi34QuV4eqRgygFxqYc8lwC9wV+6GaxNbD61+/LsZODxc54kHeqS+8Qc8JBXYwit8+RU6i
lutddlB9po7hSZ4M1sObacELb7ZQH5HjgZrBW7TrJCKyEsuQko6q1+fLontI4VBUY1GmqTEl+dU7
QSgeqwNvC6gtWzzFV3LjSyQkhoBYCoWyLAo/eeP8FVH5vmc+Mz2JQhH31PNOza30HiM/Qzmx+qkG
DY1NeN6ENzlMzE6E02m2k2+gfePegTZz+bGiNAq2zwBPEfi8TnKeZohJHUnI4RbuSbKQiv0HNA/1
VcVviBaOYZiVq8Bmu7pYh7MXCwV+YjGh7HgLdGO0arzjL3ZwfXf5BKLsXsP8ydASTWNqaHbT2H1k
kGfC9qXLyytEr/qbO58w7lo0cMGpaNHbQ9Lyjja6LzSqCGlV/Z9WjG7/m50/pZ6hB5zR52BNJRlm
GXKlvYgwbvtgMYbJlx1RzKW8NrpQQCu5OIfvbcWPppKxVLqDxw8UcUxR9X94V6KacQZF2LXIPBDl
g3pVDF9iLC8NKdhu7LTMrVdq7A3rCIjxGQ3dw1nUgEa3C55ho2LrF0vWnaRNRffFEt0XJ8hoNd4j
zhzZevh1CaZ9sTJZMfTbpKGQwSvI3whc3So/NR4qWUINgxwci2AwAt2VaQHFBx23+aplKX7+5bM7
lqveo3dygsoSJiLwURE9sjjFq196xAIZxllwLv7NmJoO0ZH8guHPRDtSwya3J9+O6BIBF4k/1JUA
g2ml6n2BLSkOIdBg+Q1gTAYTNJVmn+U9jatBnEhsXaL3ppPxEDEXUlWfGKzUdRA6xqdFNxO6qt05
BqLeKQJY0suwa5PP1EKPT9HxH5F8foFoVQwM6rauqW5kQqqjyBg7Wz5K5JQoTs/XvkVWdO3QqDSs
HQmnFgR+ungEyBS8180Bs5uaFzPcnYWB66dylIUNWQ58R0Eg6wojUXjfUgHW6worOhAgOL/Ytieq
qCcxOf4+iiTzonHt3rgPHAlgM/5P7dYJd4wS/yy/MQQkH4HIey8mmDJmUh7b6faocbaGR3BXO8zF
jqhtNGUWFuJj3A0TAXPmMbdtbw+uwGUhKJHjAL/qW0WXa0W0bByr0U56yVZCf2Zx/LmLjuzXHrGD
tvzG0FDe/hDxwEb5xtN1aSXa3ZK/6uMj1aXHcTm5WNzaFnrqayWzPFXmi1CeGwrZxMQjt/8ANbrf
Ewb37as4pjBfNyrQ5SHcxPLoQ/4bo4sot53GQB2jA6ZbIVHZ0e2ZC/UZkZdD24EqRvNEoRDFGjK2
RobqbpRiOmon12DQg5JuWJ89K3KNOud4kjEG4qTLR5Dr2de7Rr+c1J+W/4ORVvqhT+FcqQnSUtVs
vawG0hJuL/i3ehnRhjeNrB5VlYc9csRFbbEF0jU8RSQuNellN2i7VaSODUx1epjbb0zXtPOosCrR
lDcygUVAZxyi7h3Gc3At9r++glGWzEAg3ZXnkFwrFL/1DqLeb9occotFpWfvVkjbbGY1hBtxhDcx
An/jno7wph8Kyt+BDlCF0ibm4hKvH/7M2ROOasiqrVuKCTCsiN1EhA9h3crBI0Ju5ff40c+flrrQ
jd9c0DE8AoLHO3kdpSyvqgLlKEu5ozBZq/8y61qU+j+zP5qvL6R53U86eaBudHppVnGYaxhyPUAl
/Poi6xY4F261xFTgdhAY/SP5LpeqR4ypj9uIhHfYsYN20MXu0Ze6GRep8VSV/LBrPJAoO6TYr+R5
m54ao7wr91XKnxVN2IKHcxTyczptsI/glEznHSt518OjeFjPTi9j/bW44jsAhsNe42vYMCYXRHOa
EfrBt+28ZiZpW0rdydzJevOXebdSwKd97RhAhM3luPV9qTsx+16YROnvL13Lx7aNamhFQNRq7jbC
TIp7G4NvHzI69+oSsd+qpQillM2Ytk0lvfkF6QA+V2w5K4UUJ5OineupXOV31nZ7ZhI7ICsbH6fJ
+ZdvPjeBeGuJ8RHr/n76CliUf7RLzRoduWQQ8c0Hmz9l1F0VrTyUwpBlqwzkKf7qb5pWh+RHOagy
UpeygWN08fDym+Cpfxk81W+IuPRcMO7VFUXbYurgRHfUfCOK4ocinA6BDf/y/pRs8cDP5R1yY/6I
pJTt6EdtHPTJRMSO6NrAm6E2edu8oGsipO+knwbtjTz7vodvM345/sqPoMSi2Ct4vKHDVh+PHHea
iHrMfA0B17x38jl9jSjuZMsthHBGf1whzJ7T4JSdn+sz+pvkQmndRnaf1TR5ChnkWVmZPyBuZtXP
kKH8vjp1tJXc7m2cXV/ljoIIrJDC6dZWgwOL9gKhLR6gZV3kQKPCC8vjP5GV5i87aQxpxVlWbBzf
pu3pcwswAt85ujdd9SExb1zb7wLZBzyVw8Pn6dYDmV4dKdZMgZkNWqPdJFaxOkwbO1OcUi2hBfr2
c8AWJ/OsHxFiIB2XR+8cwWm6/UUYpam2O/CxVBBW5DmlbHpF17dB5qE+bbaGcQSHLym9Ix5RyiUL
RHTTIZfJUk7/93/Y2xrJCDr0iFaqL8F0FGGLlm8UXDKyJpYQJTE1KQ6FQA9qRrB6QkSN/WEsL46f
n+y5LMxfymZFyTfsYBOu/37kxIEPO0si3epyeiVz5fIgTm4Y7tu0xs0pgXAI68gpe9kTDjmOIJgI
3s5Fg9Z9pQJJIs8UNzvNqFr/YisJqpskZob2BPw+6FmYmUD9VG6AAXORwAx9fY1/B8gTDXzmwisR
mgRZQxLEFwskU2T3UvfV9kTlLVsRH9Ni1yQa+252A5UTcWnC0TkBpp0XcAAttjlLU71jCaCe8QD4
ptld1AHbaZio8QQzqqsiwbYVu9nky9z+DoARj5ga91fCFbgvkKU3QhprI0OSxs/f+T7c2nezlJRn
XRrAYVeWDIpQG/3NJ/JaUTO3RhnjkWGkl4LkU6zkKbo/GXuBQs+Ohzv4hkUqOw0NciRhdZaAjHaR
vWFhCxK8UVKwGb2brPb1oo1qCgTLtA9ZZqTLjFsYjP8DcHbvSYdDDIUWobxzhGvjEtfTRYLCKQd6
mALbef0lvirUp48l78AFFx3UuyC4XaCfRuX1i/FQQSx/VjSZrgoumGfO4iyEAdIrOWeK9HhUh6Ye
+3wm4841DOYEhExRBcYZyv4jLf+VhwUX0FeLBMm5yEqBdW18hVnUMzzY7L2LKMAVtQ+adUOe5JDL
Vkct/vBZEPhXwTRjUBnkm6fe3Ljxl5tpaRQZoN3RC3l+EQJXWnhZfrL0i4RWD1HKP9QOQF4frOQ0
Cc09PbozSH1vH8wBe3mXQsqDvUKMNBelKhIikqpgu+rDUeZO0ohhymAsxYLXuvGxq+3wVgKhPD0Q
qoxwQVMxXecCAFVmT62CFyKKiUzgWaevWT0BtxGkoKUGibSsv9hPtWUU8wTok5Lwe/NiQ9u1T4NZ
d+s0BbWe56qmryKcaP/5T/z1V/6F1msV4XyR8IFFj7C90PK6Ny0HAPRc2fPDtwO01spfcy3LhSRR
4Q3GfIrzKJc04gmauXHnPnuMOyUX3qXeUwguHhUexFPOMC2/G0EXmu0sJeav+XBxSbyJVlPm45UT
ZYToVI1cjftjBedoA9zUQZIrHvfkXLnlBoAK/bY3vmOodaFqNoK3hXipS9GKTwMSNxwkYpfyFz3+
n9OgsN1IGB8b2O493EAu9x5jB9y9dgBdyEo7KEFv/DPeyL3amdXAGwYxUrwCBDDEp54AsHyp2UIY
lK8ZnyXkHtgz+aC9B63n4kFuxU3sLKchTmYOOdDa2yJilcBI7A7u5ecmSSAO9zWepEu+WTKez4Dh
l4t301ad1/2y8uuLWx+pER1/YYMgS08cbD9B4ATL5q2rh4ap7x4fZbWJTPEaxpEtSKP3ahi6fd6S
lyvgWhaTBTJwMSilJpurWlhqaZqQ1ggLOHiyEPekH87Vftb+2yACoYVyI9++1Vl3qc2DpjSFBGHR
CXf3ZfganjCfNHlhRESLtZGR8JNzzD60Wpxh2//75li9252lSQ/HHD8xhJriIe1wtvNiU8jByIrr
M61BHLBodU8wCvGr5/ySrHZagWBe1dxXFvTMKYzimbZ2y927ejavtPcxci/KAKcL9R1f1kJGVyI1
iI97qWPkid5BOQaWFeuAFfAj2U5OawG4TqP0HK3Z8qUM7TxuAIRFG7PDFcUEd/+vOR8IWd5ekZRr
9Y7cfKaD9j+ODYuSO9v6qy//Q0CkNCFgZE0XUcsrSn+avJIC7kNMU8ARyfSquRNRUrRXHaDSxrLG
qR5ZkD1XIGFwPJ8ukE72NMZMQ6jpczVyButFK9QY6LDAkr+5wCkb8l7x1Wmvef7rWacZDArLYQJH
0CNczsXE2uJk6KFifT0J3pysJN+J/LlA9KHYHlPJFnHHDDbonhnoNZ8+Bw2GhtLGnL6aqGhe3vrI
I3N+JepFDfRaX3SFIj2VTARMQ2b8PdEyc2nNd1Eo9Qe6k2I0SXs04n0yl5uDRCcXNmmY39d2K7Ui
ECKdyxajZ12rW0V5+UDYyqQZBhZs28k5CPJMs66XHgEkYeIr8yEnPhtHX7QbB+jhBs+TmCyhC3x3
cMh5LgsI+21gNULatIOwfHLVMbd20MB+U2Gl5kDzARkqy2q4dgZVXOy3GH9bbJzDQNo4FJKuS+3E
qxjXz9vxbno5Jlj1mV8mOCTy1vFE/sBHMAfhkU7pXNO4cXRNFFbNLcAhsqrDL+lFv9Pq57zF9ggB
C6pmEYvhY+YF647+l1FLq6NTLEwmGDLztYHEgVei6pBZ39Loytp4zDJ9f3kTmI7wisuCBytfzmvz
Wcid+eWn81MiXgWupxXT5CK9isMQw38y18ViLfofuvd2+0jg0aTqjxEIgpGg7y1Gz2Ts2j7PcffO
VEH75rRF45W0pbb4P6mttTZ1Rr9nptiK9leL/+H77/8njLO+6ohf4nL2hMtUOciN5e/4O9Q6MJkm
1dIWf5R0Uq3wh9Yp/6CUSS5cjxGi23N2YxnMx34vEYNA5CVIDHwAQL3b/yioVkoZiZSfQigYEd+n
5TOr3ORwkD6xHDwOrABAik3fbJu9TIX8BBfki8hAIizSq5lsLvEFnwpUi35frP2u4pDYd9Tv6PqG
yuq4zjDXcO5z/PVlfICkg47V6uLuqt3oP4WlD/go7H5ZQ271QvOWR4W4ETyVdsbl22FRNjk01JnI
jxMYKsvIXiRe1CE4Byc1vifIZsNzvSYkhkFi0MjQwZz+V2XXI+Vgc54TT92zYP5j23tytdABQz2D
xbILX5o2NlZHzFJewEA3mT8sMSVVmiqVbfDxsX9ZV99jqvB1/2+krVc/UnFvepoM6hkGIBL5O0Z4
2/mHs9pCb8uwojTu13DYSAPyCKcR2eCxPYZ8QPs3BanitghDW3ouYyqBFJF+lHQHCwTnrwFhGZUp
VyBhGnoVBnt3yc+HWqu1NcXWCiAh5EuFmTHAHazHerEAr9Jw9tklr0Il719z9ZVYnVFJrE0gH531
eYwYhabmEg/GCHA41rNIBjIDzop+gqaUaHHutG1GG4KTt2PsNN1VCpqSeiSoc8vBOAeyzsIvboYL
bSHH3bb87qTEAzDD1wBjOH+y2dOnNO88FKe9QTobtWBcvmui3RyA79f3Z3RqdzKi8N9ZC0V+xbPB
feARlQ012MENveNCdjwlSXjuXaUEFb3isFUB+KEV8apHhO+1UKnJ//MpgQXMabKJl0/PA7Q7F/F9
BXqM9oV8hEwLaPsjGHTsQN+V/Bh+F+lmgvV1oAK1BxTku5dSWh/FXZ9pW8/l2r+ZDGW9ASLgGdHe
w/W1KKNbpE5xTCXZDGodIIqlFfdAQB7rRFITdEJmhhbYwpRn6FzZ6ILj7ePAuEG1PtDV/dRgicfd
6ssfTwB6KVaZC/uudneSN31r9QkazjN5tITHnadNCNMepa+OOEG/SjYoa3pkOr0uMGQsZu1Qgh7p
/Gbgp0YBpwbuB1zBvdeM7NwJ6UGoNM5cEKSyeaQNiII2kXlThAmxCYng3k3HdMpwemKht1opUrQv
EyxNinNhOSzzoHriDgojzXumThd7BxtWG5uZMWjsABYc+Anw/tb9368zxKIm8LU+3aLtcL4OaELh
63goSPec+JEFVwGnC/5rVuj7Z1Ml7+vgprzR9L0DL4zqITCv9W7tqejv5GqIyx3rL4oS1KM4Fys1
bcP1As10JQTESbTTnW6UIBf+fsZ5iNIap6774Xe+RsbXZY/sjz2D9oqgWyjTDqM/guA9b52SxVu1
f8aRPhVJfpQuok8vu8cT5H9wzP7nv/mxcqXe3FdIvE7hthcdY7roRw7TxuXKcPBq+vDF440Pd0Kj
ljnCYLoKTTL91wc7Aterh/P8PimRJczOAJ2gRb73gco/4Uly2EDPKysfYSrKjhfJ+P43b8Yz4K6l
n+etywhHbXrvYWXezLl+mresxSGPyyg9iaScWu6wlDjRdJt/Mtfs5jF0W5NNNz2bmTijN5ybgNdR
k8XVoW/YXwffFTwGHn6BqAkS7G/aBLsvpegZ+pYkupYf7L4KoqMoBoeFRX70o8DK5yQR6BHZT1GB
HpqnAtQuA8y3Al/p9ZUpyCP2UnJsuIC/x9h62ybXweGftyAqPiatLJh4doai572brgxNejhBfRbv
dFTIDzh9gpwdMN9BmK32OeP/f+EUn8hgWoz7zvYst90UNzX2rkVrQDkDy2dBB+be9txhEpFuzGLk
nS1ZNH7/Z3QOwEC8qFSLABgYcQNaAkeTfITofh/2YwXMU7GTT8JgLy2gtxHcA8mgkZbtAzCEBrD1
bG7xnE/XbpopnseRpTzYFmHb8GGsc+XxaxJgDZYhYaSuJ5sSwuznd7a1H9Qmujn67Ojn3tnD/i1g
rDNrqSsaj7oucJxm4f2S7BNz7kbQdCregGyGyKiYHEdXQk10f3CnWH5hh2NpJc2VW3gwT+Ah4rdj
wqtwvrhUoKRQiC3oHkIZco/0UKbwIDyRxCMbhsWahQ6ccBsQ7ZJiermW5UvVwF1KUP5K+qkg7Umt
mrhkL56NUmk0yQ+EPIC/K5oPVCItxMOwVdxK7mmSuz/E8RXg2+90C1uN3DIuAUchnRdV/nV9VggB
TW9qdhxAzJso9oyyRQ1m59Rcjv2RFBcFLz/PKX+7QPB1lQgHRff9JzNKHCJXGODqbE3Bu8l+jDPC
2zZWwHWA4R9S7A5PyOb1BMeLZqIw2KjOfFCYXrmFBvd+v9yo1u+pvwXWWbZ0YHq+Iw8IXMNkBZmN
waxtJ3f4DSSpfLWBHJGw9Q4vHWYYCCiB0g2DqcAoCjYlD4hqaWdXTE5yqICFvqTwqNIYk/nWBK3e
lmJWa1Wsrf26dF6mdQmmsADNpAh8gXPNRydJYvSQQFIEASKIBbX8T0RKN6EmMpxmbxgfMPwpnQ4E
oKRYEF0Oy1PmQ8rbbqJohRxvF4weoXUuHTAtDR7Zf5LxwKg3uasYVThZZQa2KMjnDMF+4b8y5N6Z
giMfB/N0WWw7Dlp4lPk4FX3NQPOkUK8aux9bEhsNlC6ZUvvqdsE/JBZwq64Q8UxU0MLzlYsYIZiF
m3JobAI3uRat5CGNEtwVsw2QuZY6nCeoJ8u9ryK0qAfWcA4TBYzjrKUVx2gwL4AqR2id0QjZ7fNn
rku+43Vthekx6H6eU/wS+4phdiWTbBXMocos08a29NOliSmZRq2LPiL7ScmJCTk3+LXmp8nvAgMm
3tIlE3vu/Z2mcO1MRN/TNiiwZBl4ieGL5+MH7shaYTWoq4QveXuTMgQUIEoNf3MLMZghqpAyLXI+
w7cGwSNDIPgzuIP7ko5dDm3Q/85fahpEZcIpQG4/rRDppt5Yl2swNnDRTR+4y/jqz6ViNMUq+m4o
Rd/it6Ue5/rn8sBFPxWRzUwY6fnlfiMiA313gRX4mUXlf+2YOQBnQMoyxv52iz2vXR4dB28141+M
yQ35BuBrNgEHcHSd2/0KPCyM7lzlPfys1SMtpFIR+AkdNiYFXgpFZIyAh/k36qD6NQDCROd6fvpa
W8GmYjUCj8gOaThCPk6US8NcvPv7pVYAXvcEtIRQkOM2voULR/5gT8Z1J+TvOITMVAhx2hRGpPSP
Z1SeCH1TvtAq+gqojigTWvX7llJA4D6JHZdaFlkntZUNbYtl4lVTLMSFj8wEwBIi3tKlwYDW2nEa
/CchzP9wiJOVMxVFYIxGh2nmMch0deQMSC8wGRLOR+ANzl1p4t74NODF9JBphKjJW7tj6HpxxaOc
TozhpnFzccd7H4HPWm4FiPz3JdLYa8Tasmw8agz+Zd2H5t3q1lGqCBr1bCKNTifL1DV0LuQ98REn
FrrEf7ndH+ymVKQTe0QeJRJ0hms480PpZ2NQ9fIhZrAdW0TgDUzS0k4k4UsHEUJ88XBPZyyJDYY7
6VkmTqja8zzyMPXtuSbBvEukfDPQ/do0FNc1v6DLKWY7PYrCnZk7MLjQX+r9RcOBV4Ppvw6Ub/vb
czAM1ZteOD0xwrGT1VotMa867vPx3Uxdxj3cga7Sn/N7eGiUlSQWxHxgHmRqJkj57TQ5H8Zv4CiU
RA9LL845apIssbXjN1NTrKN6XIYD9vRzR7gqRi12rHV6Y3izAbhSW4V3RhJ1kQUclgFXOXPu987d
z8BipBNmI9T9LA11arkc90tV7zSTCr2j2ZRVjp4Y6M1xYSbFY870RqFAGpwhatDZXC41ON0hEr1/
XLYjWv5pvzZGrVTezEozkqAouq6rNzkG0sUzuugayHx1IuG4jpiGdEiRwSCMSpQSt57MVCnl/agu
4+rW9BiK2QtRiGP/tFpsMh0UfXerzVkctW1sEIm60faxn3YdTCDy9MRnkr4+2dcZcbja9z+m/bxp
6v8TUmB4yR9LwpvVoNG8xZMFImA02XYdiuIdg2X9mwFMtpMddlX8zRPnugvYVuXrWondjC43fEBn
SEyvrPgGblXYCRZqHNN1jXIY8Ew8/L9fx3nrxjGtoMG8DEugKI1sZp+dWwFe5VfqiRbnXEpVQtVm
jf7ypz6XzQ37eFlv3UYOvAhakgjKLH/IMBvH9+dE4t4goCs0RnQH6BgRHrBJphX8H/A7xic5vbnv
JnR0YZuPR660PqRi+8MTNvAo28gmoXi4qwjaksl3GggV9h+nR755dPFsujpi4Lw+jyK9jgG3iCdf
7yLMJYaKkMdsPFm4pVK1RJx1HFSt2p7sryL5blMI7Bv4xSdLFWzBFUlQRjKJMZlTNW3KAdNkNVDB
DsiT2WiMwq26qTqAaGG2+SSS5919xUZTW3JE26cO09yuHBlf6HN84Gc+/uyrTCypTUV456oTWGoJ
SG7b/996Tpt9PP2LibJKzygaD8WqOu1xaQDLAcX98U6bUu5lE4BuVA5hNMVCGNyx2mO8J2yeVymU
x9yYZavk+dgVglcR/sj1vGJ/ZXX7OzHTmZn2zjq0SN0RfyXewL929GzdC7IdJpBolvp9S8yFC0qn
NWdRabRLJniGN4kOAzQyqRCaOttnwrVvGe+hFHlDlHU/5JNRhW7WWBXmXQVEdI5o1EAYk9zGMOhH
Li7dohU6rAmwhPq6d7TWBKcRFcbBgpSuY6cV/ISPl8ebT9tTkpOlYm86VZBGqhb/DlpLoYpgLyFL
poveknHSrceGLoz99Ggm+OT37pn79hML7XBbgzbgi3mV3NYh7ainD/vV6wpiTSFfSq79HfWtTshX
Tsj4bpTpdowuzvmhYnaVlVXUXKXUFYwZrZe85rz91nZYSZit9UEx5P475MDaoyX5dk92zhrYNDIr
Cfh80WCs5+UlzfZm/z73fwQi4xi4sRoa+Spu1OcBgwRaFeGIFOe6xZoGcEMCPoHN4Nds/phEsiQ2
hVKLRDvmEuXE1HflG/Qg0eda6JdwXZEDixxCUkK2UxGPa0y9q3SCVxxKTpq18si6BJgJ06dVxC0p
vOgdQdkgnhJn9FScuPp87kCWb6tRRyI/BuV4TZFmUhd5PJQbgQa/i6RW42vpcJoFXmnnz6YVd9vK
kTfYNBw1FnwWKOcehInGkxUMtBpkDLSGH/QCbteaIPEKafv5HwP3LpjKkdNvHa8VKX8l2pw1peBc
RoAXXRRtVRLcgbT/yzZtrtb/TjkHl74CBxFNcBN3RFMuir2iezueIHlmpXWeMNgeaRX31ZxEQKBA
OfyrkBgx3wTVJWmoSjpw38HItc2RMq+X/973Jd+RoChkQzofSo3DkhvAzn1GyZdTEH4aTbCZ1BUn
kVNqQmlH4ayOuhQNy7DeUpcs8rEcwdr4dAQ44VrAgBMV7EtBDjw2XtLbNlQZnClSXTThjRVtXHCL
+6j4Q1fQY9JeytMgem1mlW00OvBCttFei+HUwQxhpLTS1i3m+hHmvzEiaCFMtHga8SIzCl46rInH
syvINOdAFC38s2OJe1E7L7lnF/ccZdueMOQeVU5nzu3Zc9dTE3OfLZRH8B4KVDyWXIkbA+d3G0Vu
ZPV0Aq5EF0NxI7431zs+F4luk6xuv6hfHyglH/eQTedExS/Ue+i5AH+YRPuynNSAxtT+pFf96ItP
olnCkpNi0XHkAo/vnFpJ1gDgdbUcvo1RKbAM3UjoqTEl/wWj4vpG3DuEq6q7EqBUZrfkPwu/xkVi
28k453spk9RRCpS9cuLfaAdLpQdDGhn1Z+JR2HUw4XuAFDYAMQA5MEX6nCPu1mRXrIJJbocYSO9c
SnfYH+bh4cRucgjE+mzlb4Qv2NTB7S3UQJEiBRMS1P7uMTZWkxxNKXanscA3+FztQZA53huB+odv
Z9ohiGU2pMiD5PS18eXz/qId8wUbEhLtzvxi5Tb6w0lw/DOP6AofSzUX9ar9AsfVEXxmyULxKJHD
aYZjYcxPLscneVocMYlTdzB/AcVpe8gumX1tteoki/xpB4FsecDbAvpjKfbLMovnOI0qODqN1VDa
vhE6V+Rv9+C7Q+/sB7HwGVGxNQLAQllXSniwdj0SXxhsy19iLqaCA1YxgIPTYDdhIvUmTUoZo+YS
bYEuxajE7DTqHUVGLozAhkLyTLdQmxr/qcl8Yc0TGM5JhZxRGKIlffcyMn7ymOzONXe9laZhpFlF
g9KtDrEHBHKJ323p/nA7gHsvmd5NW5kp1xiL1Mjd5sViP6LqOO7/g+Bg/NBKM9S9i4oH8DcvEUsp
Way21EV9POnAv+TJKx4mdph6PMmTMWiNFroK5Pp6C39CZqtERWVOyFbZnHykYYMRBcosro7GKCWI
4rSTeMX0AgOcjfH9ySiu8ZNvQlZS9pzsXJNoyP6Sed5nyaR7Zot0R/oXUpLMI1TLxbQwsbYPsHOB
NjUo+DDCm491LtzgcYhQ0v6vUaLr6Z9yd4GC5oxK1IpX8PsKjTW5DiNmjkCplGquNrHUK4r4O1mY
ZvcRamflvVMZMhpNIvZZ6i3Fwj0n/tjDh4MHLtLiNCE56/S/VIoxJpeqtmFuOXZ7xLEFEF2F1Yi8
/t/QmS5gUZ1Ycmhl7TQsTQnj8RB0rJj1ECZK1h25sBO/vTyP3BHs5dxBsVWLUGc7la1AX6fvDwZf
bjYIsLn7XVmmhyruj2fKJ23m/5IUSyl6dJ+BUgNeIxnV3IuSv9egFARczahp9aoelNJ0j8aj8A+i
khAiMGWUsl0vpqN+oJu5FHe8Bf3tBAhe8WYhvXe12kEAvOzThBEyvJCDaQFdZK4cWzFW0tgu00LS
XnnnCu3C5ihpuiR6uT50PNwckbcfeh4Fo4Ha2C7mXQXwtblrRX+/d4uNo2CRXHw0vmHB0tI13S0o
AJYGJWQCMWFCxcPdAnkac9ARHAHAXYhJRt8DEXhGX8QbcESfJE3b7AlPVpbCavDg078zNXpnyeys
g+I1crWPvpY0XzWtjQd2XTOUbcmThLytjOIdTnKI1FJR2qOrStZa3wwdRLnBJPCH4pJwhFSdxUHp
3Ut2T3D5jqYC8/I8X2PpJ6hSTK3vPhhXDCYwkVepvbCKpvz9wJpbCU3Ix0p8+vAw5v2KdR+TedZX
W7sP47WEz67GrO21wpXCgNiZ5OtHSO8IcJnTrOy2N6unW+AAa1/lhNE95D6SeyWpjTerCy7899r7
RWE0SKwf685zDuST+P+GojkrjpjkI2xV4dCVXk5Yy+zE5W4hZCXpfjz/okqD8+3yeNAOg95JTPJe
3piCRZErPjeBYFuAZBdn0kxIbBoSXarMwB5+9RHqZTDZiYfWDZPHh7XNGcfx07YVhCMfROEkzM9C
teZZtjpBFGeEK1Kz8gwK+RHGdC4S3X0XkngMqIqkHFd4oTAB/8CglQb9MjrbSSYdAbsMUsTQ1p4W
g3LhJxM5UdbCNZw4q7kL8CFmz3OG4lUhFPNe0lIa/EtRxUCm3pXNdF/wUTDFdjEX3+petnSXq7bH
MMOlnlRJgovR+PDnE/N9I+EbZIB/7Ud8em19kuGzBqmmgAbWWO6O6Jh8TywFEqKIl05V+u9V75Em
mzP+bGS/xFgUF0sZliN2hfTPKEneZky1Hu1n3SDzZB5foenl7Kv5JffQT30YCX29pYTux5x0pFNa
T1lIpws95mg1WTHf4XvS07Hs3H2Jci6JRXv8vJ7jbAPpd/TtY1nsWNT1cEbq4rU0jpGm+M6TfuiF
Uduf1q09vxhaw+HSCYUebCMDuACw0arbJWkBAnTI1R1akrLIMRotaV2tfdEBwW411w6LckzgGb2V
wjc8qP04WeXkphJy0wSU/bx1eYLERGrRUNIxnOtRGQBZ/xHFOqjBRLkVNwSYTaHIIeMkKuNG4c6y
EOPve0CfotSX+7S4hPbTK0xw/RfkPDto0ZZrD7dFGpWMYfhFBjV+cK5Q1zuYIDiMUtf5VLML6eDc
5EwhcyCfQWw34RE1eSrNPaDnNmBsBgBcIQ6iJrdzxGCcS+npAsyV7IrusAR1CpjvpDbQUXNC+g51
dC28HERcxFZTBQwU+17y8bTtK4RX+Xm8rayo0NDTYkNMhkpBYFQTDRzghMpT8NoMeWZyqzw8PoLP
C6iCzzMNItokUp3i4jqw9e51eGJcDGvWH/JqYGvpWYVFopwRrW0U5OZe9Fdel16oHaP7j5b0Xa76
W0blIrLEtk+m45JuxgQCKxa/zcHrwaa5FVpH+uOJ8Zlm7t1IRU6cLpBGypnJOgp/gAQpzsUMlQMP
2DJevvB3pjO6HqzPsbodzToUwqSAUx0TTRKipUcYH9knvWtUDxFImdNr3PXm8txKET7Q7r2CXlUs
C1RxUHpp55+e/faXnx3m91z4ZMocH+VfcR3ou36B3K+nIX5pa/qZSxX/dCKoqWl1oYY2U66HvFt1
7ZhWvVBuJRPk9TjJF6OeIqIraWGVOiVauLLsE6SNkoEvNIBuLAUb5jq76KntofdJ634O2BEt3H38
zUFKk59UPeyXnDVA+URPA10A/bw/EGQM0KO3+SgGcADfObOOx8CxR88xV9WeOM2kY3OP+DkAR5pk
/1pC670ALndYHE+TEihPavXJsbs40nghNQ0q1Z4/iDngWs4XYYiQ/hasGaiihoRBvI3vWqevWo5b
mmBgPHcXryv+gugNEDQUfOtlv31aqdhneD0zxjpVeTIxeIQ6aDFh+PsDRi+M1SVeTiQHwqlxWY3k
V5lQ9cBJRoi8UTviUVZ1JmOLqxx2tfDlU4NTRpTTCK9cPRrgSWXR3QkSY0pkDNHUgweh7chyujrR
Zp42OEHQAWkRD4wG60MVriOWpYkWxobueo+ORU/Row1xBnRant43einfh+8QthwS4blUf/e0EgXS
7xd77Ia858gLYxfVgb5T4rOkV9sftw7ZF0sh6yfuIgC7mz7C4dueI9UJ1ERr74CM5/FKSt+XsftN
Ba/quVjxcFjtEaYzxigwIGz42N22/w4XXUosM/cwd/1XX49h0976vjfamxQqbOoVOlsGkd+bPeXZ
7j4TuJ49mb3Z7rc11l8dZK73cTzzKHp8vjT0jphhNSC7nW1OdH6cl2PibJyt0z5S/7KLcK5hcCrt
U9XSW3L/2qe9Atd/YQh2db1IeqESjndV+3k6/76O+/X/tod3nYazOj2cVgH7yazMi4u4JYJp0M27
4bhV/CGzkNRk+iOuYVP2/8s3gfxemgT45kRTUGf6lhT5DJpsLuWwpfShPxBBeh1JA9cbG4j4/ALr
dc996JMLuqeE1iu75j+s4YyIzBGWq3QYnEtJQ6DN0YJW0NBqKuLu5A90N3Hj4vMhznfpBg1Xat3b
hSACO6ecyG9GjywAg7z19xVFMtkQ+KrbKx0QkFVgUQMm+WY/hnWq+F7IZW51PDgoWOTzOkVf28Cb
GQUrgRhpGoNvZefbCCji9Gbv6rhbmvOaMmktnFKUv4EQkJIkn0S/2uwK+CWuqvy5XNeSRMcmwlte
t5QvjJSl5GiLvAVr+HFRxDnlEqgKjclliGBqMwTupdf7JauNWBNsHuLgsduegDL1q8uIMGwv9Q9M
YDrFqNg2TF9vUIcKgLlOWjwuoOV1QXqi2/qPCe6NQJlzTjF/XaIO91Fhb7jn2N18vzl+6oEYzNLn
EEg9TwyJ25fFRgSHhVEp4eRgsgBTdJlJpQASTbtDx2yJsiOKTba8QCH7nuaVgi7Ht9ioczB3OqTX
5MAtAJmBrDy2nYhhs+gZDhDkFYlVIayaJreyL9XARHHDVHI4iGhkaGlsKGS+Q7U5wIzIBPAW9rc/
tZunGijRSeS+zDOmfdKWqGWwDpSutzj+EQzx7iCx/2jrJzNmM4nawAf7laP2nnY+bchMjdAC5d9A
QHF8wWgRiqohaeThU6sOTsIoJBLwo5Fy1/MB+wB+2E84NI/knLZ5muZEoLyOUZqrA+XRMmbE+77n
0QRWM9Z9jONd384H46IzuwHQh+XX/TsZFyeJMrpW8069l8qs8AVVuDMbc0cHbAAl9dPtJRuOvLOD
8TglwK54k1uvOgOHa2gh1YEntgp78oMxJUNBDcG2c//TsXmq4LHxg89v8zhkG6PQzRs+C7S7L5IJ
H9TaWzEbIJChWV0R9gt5n9pBFgOAE3Nr8LpQntJYc5cdN61pRIWu/x52mOQhEFQi8oH/lIPrNSrK
IFGIIU/lDwDKEyxFSmXOsdQ/XZ//u9ELXbKC4KBH4QFYfKU90Coz3KZ2yB6S3Fng54JEb0R6OEL/
Dt6UCUTX6MkgO+EDBYrzV2tsJvztTsNIwBIpzN0hbT8+COI13qoiDrGSf8W7/iNYdb5OS1TxtcWL
Zr69JknGz9tEl8WG1BLIbiEZF5JL0FNSGwqosLcKoLJdbznt0xHbQLBqhLgOcpfxk+AlNJVhViVn
fY24sipbScdPdX0pFwNL7NmcyNqSZu0gAHOmI2UEyoVmEAgrFqmWJgQ6EretfhWoMS0LeJylxqY+
o1HdhY3vTZmY5FPhOaVcGCaffvwt86pTFH1dffX4gvkksO4ifrS4AWClsM2PzJo8zTzdRTKPMh8X
bvuWMrepOLvNRb+dZdwXqoKjXcYLFbUlDI402zSY34I7XPBL9I25WlFj1c8qsvBzSlotDz3FNMyx
3NyMofLd8PAMA7hEjLEK9ttfqeYG1fHfkFFiCbtBZm4M7vYmqqc2odz+SWx+Kz0b8tzXJrQ32tZq
qql05co7YYuFdn+gySOuBPZydFRSmwYlFPiFzdiyVpuiiaUDQ6rzu7ybNhbNiw1K5zbVjhSYoC7P
47yhXy73yprI2NwzEy08/bYipu+0blMBqwf7ELDfLQW5ybG4OPgfDa8LI0xUfMK3GjvcVO9ltUP4
kzGWxgAuwiuxlKzC3rp9+KxAusZUuRgKqrvkhSQMAL8NIlhldHspk9b3GMhLit3nLrXxS2P93LyF
1lqRvk3cXRBz6ZwFV8Q4eLkIiCSdl5Y/TZWRQkQ+5evz8/EG7EvI/gYFa+vro2JaOUJKnzR5lblP
Bq7SE55KH82IRitqy06D2opqTqLaikbV1hqFII90qImrHEy3XGuiRLbmgu0tYCfiCMxMTqfUQtWM
M9eGX2SXNQMZGtaD6xpZqbGESdwwBiqaydobRY0bOoeJkL0F28AWVFHPf5eNfqX5+N6Kk0VhNIXZ
KlhC1rVzgxI0I011srtpRjVxDAUQHjny2dQ0QCAz7RN/iXy+ZjMbdrsnhPZPzLlkKmoC1N3BFAK8
VIk/rE8W6DnYFn8FudSmDx6G3LkIJ2YI3OC6+M06yCGHYCeRLI0kI5pRoq9+g/C+ecixvoXzpF7k
L+b5E41D9Us7/WhnJiK+WkPMt0NE/Eew/LX1vHYypUTsPmFzPlic4djAR80RZN2F8lVYlJrvbTLa
fTBoyS0131Xh98RrEQpRCg60cFyPX3tPBRNVJ2dI7AMHg0K9Od46VE4MRL6kHCaxyF91WnHAEO6H
5AruWdD5uWZffszjnIzNZi4bb3LQj7cBp4SXRDnsj14Oku0WL7NUDWAbJcyUgGAyD3cgrdDacG9l
mzKAvb7wy12IVHnj4w5Im34/WUINOk5OqJtfDtUIIxJfJX61lyva78epukrka+o8Fg006t58D+aB
dspNi5IkMKYvvD3JWMEf6vdh/0M+ya3RaxkWKMH5hwDtiSNB+K1J2KIfRKPXhuzAoMfYfUUVx9rg
1EO3q6u8iOR3NkXnMG5eo3UlFXw2AtUZ9VcivxjzgYNaeGrvU4my5h1vYZGsgbj2FAO2PknLFPG0
5UshSfh9VC8rzQNWpow7NuIeJ8BBWyFFaGhv7WiMGwiGot0hnT8oNy3FgIdFVhEj+4MbiW43XHFi
yulZJFd5aVFBo9OQo+rlNMNx/1LAEv3oxjIADsMye70t+H7zSCZuC8D53eWap76DLerAZK/n88hJ
zCdM4i8honubMHSj9TSeC+srNR0JNPkd/iS/f3GknJq8vXesGIkTlPWo6evjRV5wKUbvV1XlGvai
iHoTe8T3WqnnnT8+6ak0CK9lnH37lMe+Q6rFJgqLRloePOO0z9VSmZkoHMm8xXAnsSIspSUEQC/r
6S4fdz8hg3Usomzg/r8lgaxPwoJWiOE4jwZcEBYZhQZH4pn61yyBy7WJhsuVHxveP58q066xs4Rk
vhZ1RtzPu9dJ0Ux8vAmuxgzwP9Ju+FKAF9+/9NUpKgarchQac4E5DMponHJ2XA8ZBiW+7VstCK6X
9xhbOWdyUlK4vG47q1xIGniV1b99X1v9C/HasF32Jz33+Nsec+LhNoruDBuIRowmDfHZqsCMzKKL
MAtNAMwHhv7TBNiO9LcGMP7/nKZ7ZIaTQnw4KUSfj5ZsbnMX+NvpAWk2pKZDei2/fXY3N0p33R0c
nagDqcAHfZEhOe3xQh8UceRplbdPrccpnl+Ayzp0hbX1LG5lUDVCn4N/8l1aOmrWyri0sdd+53WL
CWw763QW0J+6RSMEb5nQsRiSNsDWJPR/mVNXWhI5WK8Z4Gh7m/flp19KTg3fvTr+Ht8/4V/M7O6z
H9nzauvxmH3WNSAV341DiRztSfxTdmEIfrkvLvS6qE01+pTr2njT8qxMGfWvyrutJTe2QQ3SNBAs
lOAAmiysJnUWZh9XjnXtU8xCxQGAadNHoP3piMZbiPZJGZMLbKdPw04Tn+r9EnHqjiRIw8i2DLPb
elJNDEMXk8hOdGfMhTmfYz+quMH1Px0JprcuyMeIr1DV6aRmXzf02ywVJdmcL62WE4v/vGoEpI4X
EbQU0Qkhrt+KwMG0aKbb01SbTjjtWMoVqbDiLHQJ9a8nRiUSyDQId7v0DwNCMkR+wsUnWFXFDI6V
DMKPY3iSwwkVl+vGQrDCoguNZg2kAKCFN9NLPtrTYHVeEuuCHBxXRfUQH23m7CmL2VI6TNMTzti5
HN+HO093tQdLlibmh0haoK0vBY5BS/UZH60ttf4uETKq2gvoIpsV1sBdewM0S/oMGCHKNxfTq8SO
BJ9SSsR/Gi4cnp++BwhyhvpNGoIa647IXOQLRSpGJE/mar5DgSS1B9JFJtSq3nvrK2tj0v/KxY+S
CuFIYIujK++hm6yPJUmlkgHbeonFsNFELLIHTf+Y9rkpQHMG+SVUmAvk6PDD/1WDZNBOU1Gj41J7
yfXc7iZfeQ0/VDcDyI1C7fNSJ/9T3SQqsLp+S1q/p4hIjw8sxv7yJecfcXzH/t1y4i0kD28VUHZC
Y1E/9cCT/qboKCUaiwVtlyMpO24XCL6gKLF07TqeB2T6X1BT5keQ5LfTdqZDxdw+S5rb5uItILP2
WKO8M93o+uacRgSJNDRUpTTYTDfetdq0xRilOLD2OdzsmF/0oEFwSZSoqbSrywP19bSVKWY/mLS/
OwAfEbCKWDoJuxAd+i775aY9qs5f5deYFtF63p85sSH19DVaLBt3/onjezorwK82JM20XHob5pBE
/ll6ljCvgKj9n4IQIZ1ujrpq1aFX4VrxQwnjXt74FSrykK89cGFgEjrEGAMEedQ9ML9+1h/8DiQP
geeOZOUJyPomar2c04BzZp3BiX3d9hgj+DM+XjH/TjKJSQUePLjDaGSYkRBwqqtvo+GH2bqiC4Ke
l453q0SuKeG85W/eJn0P5IIi0FvpehOxp03HZsx8RvYLrZSUhadMMvqdPF47mFtSuxhKsb192lkM
Jozp5WTkcJ23iUiVFO1m2jLRhAxo/PRI4iEjRnA7l0CkYgOBjbQuj7pSqkJOf2d2ZSCp8Ywiys1Q
0x/CIWNF/T4J4Wbgw6FJ8QOFktjkA+nY1GYoOOEi8cRcK2+cSOas3Rxjp/tiKBwh0DwJVLIfWM9S
RgaWK5H5RzISaIfqcDw+BJAO8X6seUCEE9FgTVr3n/2s5Wh3kj8QooTaxeLb7A3BmYrTMFYb14DM
A+EZnbn5IwjTfj2/zGNg4XtfhkkpvDU2woj/3M3dpF6QcBCeZDEaHFgbX08e48NXLTE8+QQbAc36
J+cKFUt2ki868Fz1XK9OIGbmBUuy1LyktHZIRmsiREBBY2SM+PrK/jt3S/1KqX8F7xg6dXC8/u0J
wauo1ILf7VAgWNYxDe2DeGJeI+DiDTc/iB9SPynLmwondHwAqAp4B1LmebGQmVUJv+bsTxbJbc6/
8HltWQd+uPEs3ImIIZpbMy6Y8epRpUeJaBsw3dMMtgpnTtoYwqAKDpnrghEBED51cM3ymvVYWYVi
WZRGiBvT8C8Wbd+KKxyOjs+fB226rc0A44l0RBeVO6WLOjQ/KuNNo1gCPPoTKU/iSaZrR6ZaIhtf
/dgohBc/7A9baCmqqxxTfNAZtk8lM+Sc2aveb83h7r/CWn9gUUYhio6K7+Wf7otWQqDIYjO6mJsb
p2chtlMeSIOe4bZnGn/ADG3Nlq6vzgVXhxOPup8fTMJhdoAB99SzrnMKKrmJ36JOH54hzC06FFxr
ls/EEsQpJ2Hl5uas80GFDg8QxvapjcrNdoJ8pvBtsRkkYB5GiBb4QHrMsfadbFrl3880P6bAvqdN
IuZcXjgHfggp+EZDzGlCeFsLnuCzQnlnS/rv+8hHdrpmsrz1kIHtUH3KXP94akfyHe2KHCvwbi6l
xUGjRKcShTs5jvp6P4WiKru3+9BGIxm1EWjoHyPzP0+8RE47jjAVLf5MEKEF1/sdSFD9FXn/LxrC
JMKsZu+qJ4b2GmC/u0RxtT1GvKM4rpXhg037H3KiijPt2ktp8yidUbV0awAn8ELDlZi251G+//MX
t0D1dfKW0YBReWd7cyLTbWvYj/HoPLEyl5Q8juvGKn/0hmwZKASsL2ErmnqfiziBPxW5b84v0lXV
eeThouwupekKlUVO0q0h/zO07BMlc3CnGWwrRzo+mjA5tQHFSmffzpMRUK/kLPIJcK80cU1l9erK
JYK4V2Vbsv+9Bx7+aW2FOTSEfyAHghkzn1DxgiRJqNtC1WZg+jm6jj6F+FP4EIRetbwSWWMQPDfc
hD2vxt9gupb05ls5PUNV/vhoslg4aSpRsdFVI3cWEPxIOjuhcNYlaI+ze78TiDx/WRx0yCOjv/Ix
zzMREEh4SaRXtWrwbT1fH9DT0BHxuk/RktrcEXh2r8L99ZtIYwItYCy/bBliMUF6qaubvjZLT59g
R04ayZDXCi1LLIxLOm4rg5temiuyPUY1ltAqhZcb2jqBWBRfDN8XueMZWjEvTNs2dOrhxIbhghPx
axViAd/wLOsgUo+M5e17OlxIafcjNvXwtT23Ar6dEWdsnhZFwRp4sPFrcQiWld7awaNCA9EZJpAr
9bAu2OuczSyhWQRvH2tFfcOwNQPMBNO6sNdk4T4ErS+rhX+dq3xO4JKCbGoO5GMpM/LExbKpibxc
T0jZSlE0N9gmZ0vTzxMwBe7uzOaZydRCBBTN/1ssXG4cls7t/xuaQHGxMe4uIWX115msjGBP4GHa
tvL5ZvhtcYu2GqQd1RVddgMWW29sqBzzxKSjaWs5tg5jCe11RE/AuaFvSOlTkXb+H1+QimgCuKSu
A/xNHC94rdTyOmLNZ7E+88k6FjSg4D4Bo3eOTl5vydE8jG3A2HjZP4AB42uF96LLd2ZVZGvayS3/
Qu3BwQP92wdYgjbfuI436rl3WTSiGGhgIaX4bcc+JaydRQfbp0jlqweJ4H6CA+nFq8dDv/dSbXcC
X0/tywUQD/hSrkdM77dvd7ZkfDUnOuFiSFHAOCb9HP26gtSG2hfKsONBjS/YsLRPfMzWuS4yFYNt
Epxih0Bv81dhjhzU7d2ndo/oIIfXAl8kmDLS9yheDsvOXLwJ5a7ra02WusG3SGxs3t0Z8cDhLsCC
O1gqYUmMhFbGudO+QDknBAMDEAJ1qG0bPV+ktFWrazHIbsM2QCTbyOriqNytoBss2Fire2fb/gyC
jbMgHVMW0kX8d7m6o3RkTJwzDS6x44198GukYPBmGNGCOfb531wgBzVWGeuVfbQ552CwGuD0yC3J
7QhkjpRys4/F/ifV0TY31mTzZesjaZDQ2qo3jaLbAq41v9uCvAyeAcKb60B+5eNZRr1wJVsZf7Fk
YutQD2qUXcbIBfUclskfCSndqZbjqUN1NKPkTouTCnF7qPUIXVNKF3I9bLpwzYDnLj5RpdR97qcj
dqzeCyWyx5/E/9t7YqYY8lV+qvvn6TDcbuvJ0S936CpkXQm1/Cwd4zhoOCBQ84VOFdowvyOfEwQs
NDif0KQBvp7fipzuyCf5W+obaFr8xI6pwgPkLrSb9NXy3xsPiT+wlvigpbRPqqSwYsW5243HSMHU
fxeL3IhaTS/97vrYT0p9DcVq5OlerL2nOS9RAjoK8M1PwLtigdXZus18tnDTiUIl+Z/MCzAR05fG
kRrkxUGW4DisU1kdS7VDXTq9YA+BtoK1WRThRfv98UnaCdkGx1CBluqS1ogfx0QbmgX75P57vSIN
gGv/eklaesW8MOlNMOL4TUtqwL0vWFBmifpSqMW3MfY2kdmkOGzoS+lNkJygy6JMzLdMCbtu1ZMG
1b56ag6ztHML32rGDn4N4tQcj6xEh67mezevJIrKJwIsrKOvLOvvgFinbNA5lAdFK0JqVLp8j+IE
K5txUL5gw7bDbbac9ijffl893PF6zzttm1au8gS1QVmddWwgZFTarpagRPUjgF2dkZqPmUjHQh4g
YgXnqEJbjWJM64PgZ+kcW52Omjp9VL7vKRf0JVbHm49AZl5e9/3/mvA6iR4POS2nmmZH3yWzJ/D9
JT3WIMpZr/Qj02Via8Q1RTbMyLToDKAZrhYVU0oHkaBQX0biLKQ1XZYnKVVbc5FmZO7ql166Cj/G
+IvPH2bIqMK+SzJZQ2vFZxgoXzfRRcG7rw8b1YRDAz2ZCaZTSQac8TjDQ9yDyRmX7wldP+wG9UY+
zUu4cj571nQGhAOxRnJSrjubEPaXbLvzIoSicbpSDM47FMvJDGgT5MSrvNc5gUUHexoqzVKTSMqY
BywUt4662zKCPDDSV7/J7IRll+5iSpdvms9ZQLLdfdOFaXcGj9ghmP7/qLWvkmV28DiMp0NT+6z2
099Oiftnb8q+hF7ipf27xJOFM7//1e0GxDuwP1ZLXVWLEYV/tv7w+6P9mzvaocloly087uENbYZk
qmtuxZCAWdqWjEZPWEEKDxKUZvWVezdt0P2hLgKbY6Q4OZ8mMLKAo/vLNKKkMirIvyLYWuVovmeh
DduK6na/ZZzQr7/Y07bEDeAHSzeVI9cfJ3LyU+NZK8qQe5Fog8kAd48DFPdOdjI2P6oPGEDoK0Vj
hiDPHIgBCIqLZXxpwhzE+FgG1MoVRTz4mjY8i60y7kMwfp27rt2JTk25GbF6x0DRwJ75oniJQOuf
aY2/bTaU29TMbLg1MaqoHuXPLbKL9ttuQxdPBV02xZm51kllb/nYPAA0FDAKbYlNLkzUf2P5m8kO
ea3mYH+rugO5BM0r2QFD9RXBdNI2d34tOYPzTE8HkdJDbi9+DikAQE1oL63Wr2dmRgBzlu4ts8UV
J9trvtbByVyrne7TK3MILKan+b3Nic+uDr3eCXKgK8MheJ8R/r8Oe9b+weIZXivd0ML4Eqlo69PP
srNSkkRPC06NaXJxiAJg2aJqVCCHhkmxunJal6iwd5I9dyaGiunnjSMA9+CgYQpoNRKgNz5HgUDH
faU1F28OlKkrUwFXcT+lfeWY9fRiGJX5CuaQZzXZKmIBy/wiFOVfURkfgC30VQYy9XwU6ApPajZP
ywipCIWxI38xd1TpHNnLQ3mM+kmA/pTicKrdIxHzhfGgYeHoPJ1YHgOJBhSTknnzlj/oeYRDiIgh
cjjTUDrz36xv3NFJ5sv7MDxJXDzh1eoyRgI2LIwg0qc2yBABbv9+2rdBJSuD/EsJYRYPQMYzSdW+
TEjQ/AOEbcOqzL8BFT3ZLaBLefflUW3/rG7/vMQmuOdgbeyk0F4QcDxVhZ8rdpB1CfqVqdJhkFQf
R1M3fGf1cZMF3N7YLE8fnTCeUNjeMLVo7E1SFMzZgAzunPjG4t5GDXCpmDZAK7JztDHbJQgOjTO6
25byUMuxEAqZjvkJxFSAiMEd+xqA/Vj3Qe9zameaviO11uy8C3Te3FNj/m6Rn9XrW/LhAzAaayv6
fms8PTMmvJZuK1+7l5UJMrJMGDjoewq4QEPt9IM85oJomB/mjz8qg3XRrewyxOV5t4iXkUn8qa2B
CPYJGHGpfjFe9GeCsPLpw+jBmWp5Yqrcyi4uG2l2HvbrkTPCwvPJqaFFbsCCzvsInHRj1GpuF/71
bm5s4jwSXc7Q/gA57R+7X0WaCVrn7orQJmqFBDDliS9SSBdjzKEspxQPyqkZNCJx3/PPRmcUNDKx
9s8rZGa7U3/yTK0NA+sfMdP8J4rjxbxyGu9osxPU5SKhYnlfwat3cuFX3K6JaidSbqrnX6+lmMCl
UX4L1BupOL+/u99XzOtX5XTr8LIIFSq2cygzxvNP2pZzfIgt7a2uJHpwaYaOxRWklE6jV1MCQBOj
xXt9E3xdOFVSqBjvbtFqjpea8+6UbtWMwP0NE7xqQhvWJdrFal9tDs+dh9VjGa7laQ8ALTPvxh2o
8kA6mAYlYoSQZQ86sDgjj1DIqRExcfCm3sgbisI7iAUKKBpOVFIJhmmFKtk2dNrZ+m/f9FHQyS/l
ZusZhd+KcTuXGb2yV3FWurTfM/GXKUmcGOjAvDvC2P/6sQVJW16g+nKnRqXhrCzB9cAUIr/vMTNr
LXD0pCyt6rbDYpvVBJ9pOn+Pj0TP1FxxjuoGndZBF/b1UskkXG2Wzh4lFfEjHK+rX59CjuxhXVCp
wLsFH7cr3c5xcHg/u6ctaZuPd71fMixhHXHOlOIktMdDI4nlHxfgy+MjSmdsfgXOAyhy1zisd9sE
wD2ntHreTtgHs/yD/nGBWFn0J4CCldbVW7N11hmYIfA42nzw4E07I6jxPee1vc2dZU14bgTFZPff
OYf3+5FintBLXgASzCUpvtU25NYB0zOy5G8i+ozzTD3xMysKdiVMi3EOUh6quvc4g6wCKtk36BiU
IV2pFHSApxPCer1aPNWoDrv0CRn8abkvjuFteyZlpKu7CFCJ7PA95eUcvX+LZahiLw7PjQIUmVqe
EPUV3/7h1brqUMMcbv2TZXz4roRoTMVvwpMLa0ry4uOlPq691isIJrKUhgjugkAsWCj6sSxs8ZL9
8T/F634jz4Z6gOTDc4vEQwVDsMQOj7te4+JIAkyoqggrqIFBL6oBAkxYDNcgfUmNEEQtDytg2BTu
+kitmTJ4OrPCvG01tKsDhENPfh9fjkWd6vyyK4g0DeQipgZGvVs9+DgdKDSmLzknSXgzsh4rQfKe
iQ35RNs9cyF8veaKnRUkBMspdG744pZwYEx00MOJwBEBRo8cKyw4d/TEczklqbEk6JAwMIFF37SM
FaCSuX3umfDks7teyc/dHlkGdhRirGhcYDGw901crzaEG9F3WE+c5B50dEwZOIgEQzJeHjQvlshw
3jNHBED1CNBAt8jDkydekyZWSiqIkQaQbcDXkesuMbab6g3ywyMqQyIg37ZmyWjKdE9BURxBF0zH
ut04Gg8us40RksWiCo8mpyxOVvkzfUkjWl4M5Z28RiTibn6XZVunuVaSntbU9tS5IXBncrBIhG7e
sb+Mv7/kqv8rRYM8HGUVwN0PWMLrEQ6tBz5RUBSqqx2iltjFJISbyK3V8m48X9x/fXF6u6EKjJym
LayqDKct9zBdOEQRNZtaDeFnk58xRjrFjEONpJmriJY/Xxn3TQ8uWFMsIjB4qSB1e9GFzKQLAd+Z
30IC4nHVIsh48GTN7R4QBC8AgINbw163Y4gU9GI0UMLAeedUfdRWUgLuU0CnHF15/vollWS3Og7U
IIc2kyqDttXnLMvcJqyXz7D1dBSXVl71T/jRJuaduJ22AOdjQKsWKXAP54fYjvyIbNGPm8Dkb4Up
6QOfnSwhwb0jNV3qGruSobeavaOSnBHpYtgCd4vBlznMLufZrNMAYD/+ZMN2tYucgkvBGlprXeC4
+sMjhI4oiiMY7zw7BKX4tBEEL+t7BLAhhUx+BBYoXc//NT/t8/F3MB7wQLSbLT1PSdNptbkxbO4a
mRcBrs9XhwAspiNh3yCCgMwDbM/uQOonP952u7iyUfHdK/hmDXwRXUMuygg1XJbdIcfsyH8X3GGL
0YcxkluikdfcYQN8SwCZzN8DRVhfL56PXl9ZYHKRbE1OQ0ya6tiQlSnXuFtjKZrRSHFjTTl/z4UX
XeAJXrkZFpRRCALa3LT6nKYy0zXB1Lj+Z5jBc4ImTlW14txSw90Fn7M45KbKY34g5HDTYDYxCzPJ
fRNaaSMSxKbtYjr2c72Vlu1ugOaFOZiEnWVnjlEvUHtkiwv5+Di/SoLd3f20oRdpj744gl8fnznJ
yHy7BGLtGvWvMYf7dlNTAxVR9HgQuvSEB+gGR3vB5pUZ0QhK7GksMk9i1p1kJkTbUkuD0dBTe/T/
csyCi/9Efcn3SGq5pX0lbSXfbDp7S15PDAu+QJW8HZwMnHlJhwz94/IBJGrz7RXbAYFNHaU70/jO
zT9maB2bn/DFLQIpmjnd9tQVRwj+5lJzLsgTN1Tg1RSuuaPZaDWh4CSNIPc2Zi/h0eFkYXEEbtkG
aKp4GfyH6yWFzF8D+JUgvDTSjDwyHClbVBZ4GGu4ruMz6EWv70M2ud4QjTWI9zvGhMBb02MPyG++
Hmw2Rr3B7D5r720N71Lh1gxDyKKZfZylaZaalLnphevYw/AUZPWQPF7Ja63rSldiCsJI36DKwPAr
Zfdyl21V2KzmTCjxf6O/N24AY7CUJSru4cIBdo/nGCgnI30XrGrGzg3X0hL3sWMDuiJU0A7cu2la
Zf+g1NkDTweutH+ogDUphUbrnOGJoyZoQ54hBWrNC3DtMfTomgXaKSOqy2lpAsYdoRKnlD1381so
jhyNlwaU2X9KQbsISAetg6Y1VTSMBxokaB0uyI9niejYKFc/HjZ5h9KKw6iVr2/e2mrjwRhjiW+t
z/PVQRjYsHS7LYLJ9yLjjtrvcESaNj3bo+6FSBzhCgR8807OZBsdxWcbUAt5Vr+SoqZu8VKBPw/I
0hFKI4z+b3PGu2Xmy4WSccY/Gb2lb0yGbGcXRNPu4It/lFKp8BeRqj4xwl7iVkVGDNwrvtvKmj3o
cC7VmWbHl2tBZ6DQ637WqKLQm86gt1cWZSbo2HxWHjtsRLLvSAv2tjo3162IITHOrzEp8o07ffVs
VIKVwzhlz3ARd+/S6unzaS3QPviUB7odaHNYF2uXT/QrqYSYbdMG2qxHpgsn6xpO5LkFGzLCxPWs
V/LY3KzfZO3QfrvYEt6d8txn8f3nmgK2ox+XZnYh1IpMzzWqv5dnai4mJRd50bPO9sC6WO+mBGYT
WbW/oxV1tYI/2Yoj4Xvw5ZPlQ7GBL267uU0GKIb7bSx7fHGw7wndE9tbv2YZ0e0Z+tV0mDbfGQfj
GORL/Kqgs5lf03v3nXLl5VI6gGsJm2Hng9XAd5zTDW0vr4IgWeFk6FAKmAuJMKnNeQC8P+JTWc3D
TtQHQ3XCWteUzmfthZ+VJpkTZ43/0d38CqTKlN7mZcSDGdSY4gzOJA6cTT+mSu3uYgTB2Shj1H+y
xQPSU74YN1NOuMTKkfASZmEPSURK1T0VSgjZGOXQul+DXoS06n3KoY2db88ZujJ5xNcDPxFHRYoN
57B/FOC0QoDol/PCqaslz2iXvt1X1wMI8DxkYUxJHX/NaS8UYGHuJwmyiWGcinZTrMWAV4zIsxqL
Ymb6creOyz7DoMBgklu2TQq+9x04tn4TF98iQDIGtDxYe9LUxnHLpL6ZmtYMd6haZZoPW25uypZt
UzUzwK61FpVu+LfXXPMy8Ejcaq8gDQ6dr70l/h9MVKUKMQX97gROyUjcwZ+BWuOg5/JOsYrzYomM
SwNlY2Iq+P5cD+YoSnw24sfYqCMvzOj47ByNr984OdxwjUZG/vsKmZj0DoTPtWkxnNxF26AEhnW4
Ov2dtvAhahTHju7dyz9OZ9wW9GB9PT6QEG7WP5iU8hlB51+7yoWiurPoSRy1GPd98GF5/ooMig/B
hlWcIYywtibiyLviT/4FXyrBH5gQYqgzXRvy+lwdhrDC3ch+RpunaAoawMWSmVKR1rgD8SBj33el
h3XoGC+v/c111AQ5q7HuI9EjgW3cyCK0KztL1JMqDO98LstJdZCJVmdXtf8KOGbXcjEaUKisyjni
dRQ3vx6zH95N85HSEa3EXfMkxJ7F2c9rX3O0shR743zGj6/4rIlM8xgJK3/JFDQcRi8a7uFY5Amc
PCzFaOg4w4AfQDR3DoH0H19CEVwhdLrn3FSZoCdQ81BYQzk9Wfahv+BSWkQJ0vEN8fPfmOvqrC5O
9Un4rtrl2Ie1OckK1E9NhckMe9XpsDtWKABr55phm34QIE6h6qExpSv6aQfHlr3RrF4Hlz2dIMdL
sBudEYmj2fV+mJUz05JerzihNRsTBKDCGSe84jjF9wefjWz/1qQCr0dfnkMxlvjW7qGSCTv6ogtM
nJDJ4Zc5Gl1TAYvoES5CJZB2XM7YtVzPASvC+KDbwYpdCvwc+ju1YSaJnTLem1JSgXPeF1NYoVDu
q1x8Zle1MBMTeegK48ALH70Itbv1BaZ4hHIh1nnBsg+XswCVn/LqJ2rI9gm/kUDC5by6KFGn2bcQ
G877LCj7gncuWW6dpUBmNYwVb764gqVNSJ+mWJQmIKfV6+eYXUdzhl7kZiz31eS2JK/SfSSlZTob
yO1K7zB/jRPH45C2D5eM60CQXRF8fi9D17VA+UWvMcPFJX/rI4ek4gDAMLXjs4S4W3h4cbbBWGNs
4v9fTl1oKbQ6WXTCyU1F1JllCn4tiUaNcWmLds7UuSKHs7Yc+6SujeVcmBR/SEtqhGkXc+/uvNuI
F5m7TwDulqeOgUfR8G47LsP1KJ68nlMHlu4KfKERMa/2WZjS3VkfJn85igMavNKkVrd7kRZknucj
V4kgIFfVby9dZ5Gcc5YuXOiP+Sigm6QrS46RpR/MvS+YGaof1DgPSCY8w1wNLJmBBItjD2kr2xhW
NaOjH/t/cmbgilukIUcRFCjHIi+CNxrCi1iX4pvQfU59ji11vcgdPQDikxnmD+Xdp8Cxzbk4OkV1
BH1pmRvRZapOZQkoFCMeBAT5azq6OY7nfGU0hh3LNGoWv/uyB+ZDbuMQQYj6qdVcylU+lhIHeeza
w9s7LzcgZogkCPtBd93mWBin0kR41e3/08crC876rN92VgFVQNdKLSOzPKbO8E0JCOpixR1UaNzw
MP2FuPl8OEr3aZA/SqpvNWJbq1x6uyN68Y77/OHFqAO9nCbP3dcHA176RSvQ5ZZ18um4qquAmncL
XNVQEt6MoPbaghPc6tkZFQtr0ftnBRQQ2tToYGgR92ebYpFu/QMznxTnditocFHfOHSQXJ/bOqD1
TIdUg3EnsGQUArryHoPjkJIX3nEr+1bGztRET6WstzvRYBlF7C3/iRt9Dsd9bsgszw6pMYl5dqYP
bypRmXn99pibef3IOXSHypMZcc4N4IkXk5jPHC/yg32ll/KVpIjVBx5qkzwFv2nHQzIbeHGqi41L
fMZwquetKrv66Dg5URIgxMhK2jbwuhpEe/PdnpgsZEwt9ue/HbSjadelcEPsz7lYyHfF1PxzMwiz
EqSZVizlivJe4xPHP1PXdVp5h0QAWmp3P5XzPlrhGdHD3nm+lbq2o6bSE9JJdXfFtrnurjM1CTtk
bmQB2hW3o7ssGXF7HIc+hQvOiTx6XqlY7/V3Z8hGLZXMOOp5PSUHnekSJcgMXgOIy9LnCa9tWQhI
s0rYzLwVG28Yw6sT1EywhiUMUGhKTzZJG7W0f3l5WiwjnVOmBavBK5vRkTA/ccGw4RQ0FzYutUdl
97jotJjEIhZDv1tiY9L2aif/gJflBgupoiM0POZkaJRo3mp+RZ6FMwEX5DuRevwFyodQ5Q8YBD4m
3ZvGPNt2VstPIxIzCwOk2LYduyNMgB0KuyblR2lTSiwQ4xZwAq37HrYiB4lleii6EchaSoSai6wX
TRrzFZ9ECkVM9AFywI11MIpjMkv23zVE0bAg0m+h7nvRpBpGPiQ7anqUR1auGJQD38iP2gX0WH2v
8yJa55zEC1bnMrSo9RJ3kmkFE+QuLLrm2vmmELXydPG+F0dGs51rYmda5j2MdFi3xJEHN7jaZm/w
I74nk7VuYEUHymqgybzelO5qFFbs+eZFUroUdrrg3ZHC8IXPw6acdZFZDFWgjETvRZmha6yZ4aTO
iGP5EnePdI/KCYgBmQpBxDtdSXfh1FW/Dnmyq53I+e1bYpICHUnWf00Q0/A+5wuEHfBh2w/H7mjI
hkv9GfmKPdAofNA+mEYvw0CQZijp4RTrrCACD2xW7n9awoCnhXkGG7btgh4Cvl4WdhGQBP8V9NCO
4QMSeVbIkiMo4YvuHDiaWZfuT0Nes/sOVgwLHDNx1qWIVVlhgRjRVw0UpgRuN9LpYlXND9MqLElA
H8eoNDWrUc+Sg+NVXda7iFms0oyyH9HEHxOfIPl/g07/7QQ5JJrxiwPNUYmFnORClujGjNqSpjLC
/mPLECQAR7LsqSlFn4sUN29r4alHuVmvVZ6+40qIY3HMavvG7IMtKxlgIKFxfl1id7j3QFYVn9UD
omJJBqegoSWYMfH/CuVkLkCpVwkGAGNfnRj+BL6r4rA/xPtz5H3iTi18j/J9B6CZdtqen96Iq3yO
goiTmPgz/y2LHIYzG/zX9bD/ZMZMhjQtZYVP/PHeSOUCtWLYEhCysJx/Y+VyHR5JBv3zISGzglRB
KxwJah1lKQmNI9beT+Y+xtCU53saPdpLVN6CP01EF7Dc6m2y1K+1YJP4p8hmUSRJtPTU9kGHNXHw
mXWLVDpH6p/n92Mn1OyMcyCL3cXkMwqOkp0ZtpisEfVMcaoiEJB4Qt4lmz/eTE/uZhDksFwrw1ME
xa90j8w2B230ZbJ7CaLBDYyzmGXRkw7KxyHk47ggFpuIJ7WXM+6XfsKF9qcDUTPKerR7lSEO2f8W
ETtaAkABVCq1uyIs9+SmgdFTdnbl08O3NG6tbBtT9QjigVtgO92TbSIW6s+ihq9ewk84uvMYgOEW
ecNo78LxQ8e+iygdltCPvJ6ffnEAtq2ZuYoq+Do756LOIkhutkCCz5NQq2ykWpJp7vG8Fqy+8vSJ
6R96+4g1yNNhAnMWk718XSEu3BSmyHBXNGqeY7RK3MbiZzGk5Lk38YjiXuF3oYne9bbuPip7+FwQ
yPXx/eDh7uc6L2PZDEiHRtLp0JYvW2tCKc14OYuyTyPl2PPfVY9cJ45lpXXEJvql1Jh3LMQUu7vc
7AsFLH7Q24vqmAqCTilSY3q9oWJbFiEkXAsathd+3GuHMhsm0l46hAQ0dIm/K2ZGQPG7Er+6lxgm
x/zoLk7FfXJ44NzaEZWjk8SAgpXndoWK6JsEh1RiX/dNwhcpXNOtS1Ieqz8ZwvZTPIyZGQrUebAu
j8Tr4Sybpb/Tu5LIGTBvo9LOTcrFq5jwmpjSwkNmGCxYi2Xn81NDV2ZS8AHSaNRBwVoy4iqJTeKP
QjAirauA7n6jzPQz2AkLNLFxyMIjs7eFmy5KWQFgwltoBlazLwDIIMTwgZ/k+LhdqDcgIKyhcPXZ
T9V9hfC2uDzAGPEJuahl0+PcIugLjlLz/o6VbwddFM78wPDSx+bOYSMKi3FY5nzhLgGMPqmRTmPt
JhUBHs2EZPtgz3dmDndEcgXOnUPY5euIZRpr9ObMDPgKMA7qXLSGCHDMWNnwJN8y4jCBDYvKC2/x
3en8CIP4PqtsCyZTmN1pXomDlb65El+LkOIH5lmj5QkuUtdsIBBd+i+4XYP32y217V9CZnNkTdZt
bNybGB6S+bQVgSK5feVuJ2vl3+mF7zOO4rM9VgSLpmt6A4i6PPL3z2rj9J1GjAVVOqGzFvYqMF7E
iwgAx7SS41CLMTS1/Qy/IC9taNdwsuiBVJf8FkwipOeFGRgJpdhsGuzbb5TQ+091KUUOC3/lr1zz
nQnICHUY8++97m6OgNuE99ySIorhN6htuGn3AV2O6O9Bpn55mDX5tNROwNUTh1MylebNBnigsNgy
AMVg6fx08jten1RNObQAnpMEEuyTed2VRBlzZhz96AGqWR1GQYk49IcFsJtW1gCp6rcMY9RqPhu7
lpC7fd1zgYPzpQQr+a3e29hsfQgAF/eSn8oXfrgCKMa3VOodAQWoX5QvkJ11GL7fgdUObC+9SnXR
luZZFaNYla0a37915riDf9dpn1A8CjNdoN775+LSypPAfJbkmCWh/bm4kCAZq5q4+f2izaKA0+vZ
ZtS4sQIVYRrSXbhqDXPM5533aaUvl8mG/hodbmpgZNE+8NzO5IuCj/PmY4ImbtSouZpFV+FigDz6
y62Wvp+QpS1u1fEbmTUf0N+EjU5TeT2fL+xdUOyBvyYSw2v8I+WTUJaOGYA7yZSA1LNGimHqCn40
ErHRjg9JpGn7445DdRFQAWqIV1fPWCkRhe7OqH9JBhkySR8xzJWFMZHoXDYZwTG29j1IT9WxStuV
4BF3RTqEfuHdbRYAl8mTEtpN0zg8ix//N0YIaICf6dO9bckG1vXVHaSUcEGzTmGaGP4P9ulr5Is9
VUHZFYhVhkwSCVOwEOOMi/QRR0FjDF0GvgeJuHoslB0JqNNEjW5hOFYaj/w5fda7QoMDb9oWg5PK
ZIK5Vhu+EbOPXR0SvKDOr+u3EcuO9hkkXdKouiOkB/KpkNYvLYoNhQi6MEOpvqeQS2Q0cL90gGbx
6jMUViYnYhmoDo++yFIrHEayzdk+3ffIneGwMFCrvDW1wN9F7rSSK+xSNRBb1btRyeSkECEq3ffc
MZ2YfmoEQQw3kbjR8wce2GJ4yW9kJrka354XDFKs9RLcbS/G+KeWdrhJy+JVNoBa7lTUU6QF7PPK
BC4He4zlDwxRHmfNDASrKom7G1s5M8OQNRZg3qy69dIpUVINgLfBh/usPz9vczfxdITArxscU98K
WWRH3iOvsvsi50yp7lZgc5BGbIA4bVR4DtvyuocAuRLDvQoo4TUaVVFbty0Srn9Kwfs9PW7UMAR9
DbkNuvFYmatgXFxQ+i/5EtXMPCOUKTzBiMKZ7Y+/ZMIjTioNv6eRtLIGqNrwD7+kF9vQ0ibuN0dM
snXejkMMULB3LG++ug+uDFwtwL1nwrWGHB8KhjZkESc9ff/mtL8dkBFyXjlNkbWI3goM/AmAD1+g
TL5ufP47//DOywhmJS3rhkc/SkZ4CogGzg5hM/2kmR+NofU4cAi4EDP/pTqOvg7BfFV7pETt5Uw0
ssXUYNVr8H+KE4t8mXt7CRxNJmwELwfj1ccRNf3oE9YYglhGdUZbz+HvkQCjFoXSf1v8gD6W6+wv
zwuGIlKtLWzGtkplGibw8GVjhSX/0Q3L6zhOgyjtWMkURaW7CciemZi5byanxNzIj3uoKu3G5JBU
asNIE9n+j8ZwHGATjJ6gYqBdVLrUDcr+Kzr5lBY7993fK49RqsQohMfV0fBNM7DU6PdJy7PDlssH
U7edHRdppDsJOVTkmJi7hT9ZwL7iw3GE/fXP5QS/oWC54t+5S+57aMbZbpBNfXf2UmlEDHzMnxdt
/uYqRtj0TMgmoByjsx6mmJsMzDZWIhFMnpAtYtwQEGqrXOwk+u1vYYlLx+OtBe8ou3+zWPi21Kyp
CKRUagMfdUDlGpO/Nii3l2ZEPl1NRRclS0I9vxABJ+Okvg5F8V36HfkOggcpmyVD7BQrGy1ydttH
rhQzO40O/lKjMoQIU0W8u+gKi5/WU5rtJtne0B+YDfWFuzx+Vaj9V+f0iOPBhxXpZ+13nWeJf1RK
fJL4ph1gqMfhe5tbtjy+UnF4UqYwd9k8v83u0SexEHwa8VFvU+RAhPYHjzmnrOy9R8D/Fbq6PRHi
zQoNrDgT9S4e2SxxJ6WglmkoBi8R9OQERwjxgOp+9St9+3xRQiepyXgLYArknT5zhm8xFvs+oYi5
yfcG8UzAwGqhRi/pitHbVH0cIY+kueXOIHJfY95RNgasPYHUFu7y2bm+poSgIEZQzDcO5dVhiurF
nVk4qXaYaJ0/9NkublAlD2mNyKD3hxxRa0YiFdOC1eCqnjRAq93gJrjLIakDxaqUCXSubDp9a4LL
JLsIQYoE8YU9A7LC/WKh+XRYmPntB0Hc6RRzn+huklojl6YlEUSXlNkuE4iY90e5sCaaN19gO/TK
T6O0mCEYmetQhZ8AJpb0yX7XWbeU0QdnniKR01EsZJCIq0/HCxLP16L3AfTgo0eUjfKSCi7ochXy
hHScVeIBoprdtuah8iBQZxW/3udZzP7KESXpPnCeZAjrHum9MTP3qbvTZ9GdtHZ+jFqExWQtroxT
WdjDmdE7lqAqXqj5fmzFFFqQwsrxSJy1tQYMlJA6/2EkT10t9veCStEYIn4Ca9p/LM2qQOs2fX1A
C+Bu831I01E9ZjpEi10Ny+edg/cEizd+5YD3mUU/ree5mI9SgZkEJTzHepq68oa1shpCdVR5Ehk0
7ezernnBZiBkfcmnQTA6H/USGm3e0ZIB7gy7RpHJb/zFv55k1uvT2ekMajrbWhR+XVNMAvhma1k+
bxv3jprEWqqd6sPJSETbIrqBy5mqfKn1KSgSPnf91LUPRWFJEi7UZugKVNs9PS+dG/SjKdz0kxIS
EU/eyS6WBPbrln5W6YsfwF0/Vm2d8Bj9qx48JaKKtSLdyLflsc6+tnz/Zy1layoXlyQCNGIueXfH
HTJSEzqWk23cREKZe/VYG1DeVua+IhrXHYeLonUTdlDWGLAqW4gp/qlKyCZ/GfdEmRTQYvLfRj4V
p1iCs0K9s0AhUBZN5UryDK6R+JvUPZn35rLrxeXJcCJ2XxWCxew7WpYFY47xIuIHJ+dp9tppxFhX
AkfFxFZLFfE34wGSLIa36C6lGYuF1Jg/BueD6h+DQYdCA6b7XjNUZS1lLrM8gzmBH9W/QHKuWTh/
CXfuH/ggHLM9E1AbiYNkYl/ET5IX6WIwbduv0+g6KGEUN8nKrbd3/ZacDve9lETbzsIUzTwDi2qu
IrRAv4m98D3aSToDOLQS36RSuji2FlRCycKml6b+M93u8IEBzaYi8WpzeB+Gak7DpnvSfRbfDnE0
t+D9BdTBBeOIOxXUT+0tUgOJlj5KIynd5bLY8s+acaxZ2l8fFO6oEE6B+xCv5UJFSgsnG66RDDTf
5EWUqIN+EhS0tG43oq0igGF/rGjrCYS2nc+uOlMITIDeuPMeXVqYkln5sOtk2QAsln79m6Hf70Tn
Pu8RMJhAIyuca60azNeNZfZnH/GAd5//aXhgrHXeSyOb3V9nyyIzStA3qnQ9mxP9fdZZ0/KorfwE
Cmb0l/Dsq7MmpbjIEN9whQQBih8emn9eoR0nb7aM0eJwSlG7dwxA7usEspL7Ou0WqYS2IxufHJvV
dEA8mD10RdW8mstXQWuUcqG6xmye+qQTX3xTcdMB+1K+PnOpnqXA5axzb6gXHvAHnZAxZtWj7rtK
wOy+YxYfmyxQqaMyiP7r9VTijQuIQtp9SQUNjA9jz4EKH/+865qovSmK56pvvbCJdD2EcI8ErtPt
JQoa9RCjs/MP7zMuIh4hwqmU+rI++yIBisYqbbtGqiZGKJHLuNhqVPwYJ8p9FqgbTo7A1UkdEnOv
77E3jSXBIIBtZsifZfVTX1D2In2SWsdPujsCpEen/jWlY7EjIR4QnCdFrz1Jws4VgIO2vNkok55B
+uonwfRjHEms5Uk6S025snoJ9Qy6px+jrYRCynZ6FvX3CSfa2twgQno7VvjlnPtZsjzmsz+U1tF/
eblqFwM3NLgc8RGeayoc6eTh5ZMqN0XFzZ/K33NvvbVFsA/C9j/ZZ2iDWO4lmlzjcvtJPWI52LiE
Bt0FdDB0O+gIzaSHcWXP8PDbRKQGzQizkpqCZXjp4nD7njM9n7q5UIm2FOt1RNY4daHQ7xsPuQHD
CTC/XBx4NShEh/SeLe0ASMjmrNi9MwJmNPh16JTZUsMPvYmj+nBJXU8sJ7nbXgrmf82oE55cu99G
ARZ0y1pLBmAypdkVwKVDuLQFf+tkuek+Wjnk59lsmmaAZrPYcu8VHanR/BpmWse8ULrQzHHP/B8J
Orq8wbhZ6CDG4yl84eKoe/vSCfTL9/l2YqvwUw/YsWdeXznlqxaQF1b3C1YgmrakHcimNIBujhLA
XO9+Z0V6AAE+jBCKpH9KiCY23p/0BRw0NGJFcZKtwf6DffwG6SAmsrExrqIPsx3kgWhDk9Xor/H4
sa8FKqPUS0EyJdzn9xprg44xMlP15geG19BVZl+sVuPXZ2OlcMtxc6lKnQd1mJe5ZgBuFnhsUAHT
X0BxdYB6jbXvo5XtVVwackvtIAqTC6sUUHZhYUp/fmBOI8Ph5yifCfboX0Byx1dIrKvj6fUk+pJF
AnQoSj0ZuP9cX72nxOmaxX9nJ0OfuStaamZUZeKnO4F7XQ9L1ArHvMLqMO0U1PXj+K8ieVv2cU7J
eiPwGyPeD67st1SylW3MmsIB2smr/tSDf0PNRldt5ZcB2SpsxoKzHZjGA76Ei5cZ8/MXpHwibhKo
QfainEV5Spa8t11RAcBrNFiso5sze6ajkh//HXrxeTfkgKo9Ldkr/LxH1UhiSpmr5v1gJWx9moMW
2hISxYYrPrT49YYa+0Nyjrg0FxuayvRRgrBHjo/m521nSFVVupuP/jTGhgrsOs7v8QtJNLWHWYZ1
QFwMC5CX1XnxYTQzlrh4yMlns4qRSpiodAuGzgq4j6AegEZjj01ptCUBoW7KkwnzFkI/t66fogCG
GUuIX/JVv/uvow+ZxlEp6WHpe3WRP626e1Q0c7y+BrhpDZgpfce7+gOlIL1hkxmaewPVvhfgRlZv
fBkV6W7LDhC2XAijvJUkoFw4uEiqOK3T5w3vGBg2JPaUIlW6SXXgfRTSxdX1wkxSGR/u7KVHkKUd
Zrrifohd003zG7fGgu1i8NZvq0zhQIudRHZnMAXJg6wm+JDV7bXXJ7ADmWGnmLOXDf4WQ0G0A0Jy
+UAenzE6YmuqB11B5wvb8Myxqo89heVlI93Wje4X9Vnqv4mFVzoBB4kS67k08qQXt/uWdHkbQtpX
JYkSelt0fJIf94rZIjAjAqEHHZbhYLTM0PJMTUQrYsYG8kAm+HbowY75pc4IYtl3/938UFe/ISVC
MVnjol/EuTUK9+/XKmhUkXUDpN2MKgvc0xi48alDGx9SY/xMSoHcuy08vJBqe+Sxti8dYadrcrIV
lo2kQstpyjkvHVNZiPlKICns5Nu6H39ZzGHrex8ad6AQ4m1lIy0KcO+RSf4sDMRt4hcv4Fo+WYOg
4MWOkzy6CutmXyi42PYmqgQHy9vIRIrDw3hk09W2V8tqtRQFTdwx39S9iYt5DNUtq5ZEJ2GSG8yp
QU5K1HM/CgPAoY6j7pDlQKIdERGVhSMZnNQwkqk4Rubefw5mAUITaBLrMYGQYfuxAg95wUwP1O8t
onlRtvkUeNi6lrON96/a/uMC1X1T8RZSNCz+AGtSEddqiwRRkPS626sXFmPh7n7G5TGgiuxptf1B
KJgUBYsx8F5N5ZKkjgMyAWds8xTauUbywHsa+6TYF0zui5sCuxsCk6c1y3xWCP69absqKO/EAFGu
+whbMKqkbmB0cq3/SRZUe0RyJOM1qZnPi9a4IYY+ql29XCKJNWoHUPxCMdY8kbIqH2g1vXa7KVE/
IFMcS8aanSQowU+q+tZuUOx6vD2WQ2ou61u0LXMedz+6xMZ4wO0MdY7sXvxeS5o07AnxP5TzDRuW
SIAPkKkGvYvOvkdM+/Bl7S2cuPcyuwARBrmzMfSoPPUcXb+vjG2tdpzNE8ydNraRDfIZc27XksoL
M2MB4Q0jKJZpkB9uJmV/YwIDouSijXDzeqVoPAAZUFXOmAyrVO0xUIigUgLLYIt/vZ9uXHO8ac/M
zBr07FsKktiGXi8y8a1N8HeMFRAsDGfkUgZIUoZou+2/3UQnCfGkt/XAYLczGRS0z8PAb5zd1fbK
nwyYTCqnUAiUdEVoOhPQW/exYbTayPmI2EZ1a8cdlMITUUGhrSKXxciAp0ux9a8flJfMlUKc3XUN
sIVmL5OZ1bGgaLiLOYfUVnV2aF7RFuc8xRdI1mnliy7Q0tDg5AHp6x+PVJqEndjRLCYj89MxduyW
GWx4s8rKNUjMHe6hSg7m8SE8454tVZEEA8rDp4j1QybOeB6qXlRBdY6r3TnYfcYjhcgGmUD3sPei
+FJBot7zQbWyT+Nv+bRmMK/OUylzaxoXpo0VPsvHtLhBH1gIMrvbSBrtodck65Bqhae3TJ/M/xis
5i/SD9JexyHuJQILV1Q0Kru79khbUZzf0T300j5dd4yvO8LihdKvs4BnS8GTDhBhugFhkbVkMc9E
eYuw2NhWJ5K8CvdTIHT61U/w3Ke2AuP31Dyk/8GZtMNuIREKvKuv5n0vKYNZkN+8G7Jad6fnMEZ/
C5yIf3SzI1lTBdkzBNRLaC9O3GLPBv7Hys1t0qY42SyY39gm593C7HL/JOo75MWnHA6WpkwY5liG
J7YaiIgTR6QUnM/Anj9oV9RjQXUJo9bEEiFA6SMqQ/TmAn36XNz9/z4Bh0iqzrYltiWJJMAIFi+h
dWvEt9EXBgCUnJFTvOCbNnnc2sGdkibtYvjOuafxZwOvp52iOLGlSTq+FXgfLOat87yQAFNzHmmU
HrIh0gySC4jmprSbF3tLN4RntOxSaJ+jTsGNs6a35rKZact435By8glHHsmPhPi3YBZRIGRdI1Kz
1hYdZC4Dz0f8tAsmuM/vJyxq1mv8y79xL7CaA4f2bIke079Pp/UzM7t7RclRC1J4wIUoduUrhflO
QLaLQuKYPYRU1v7FAiuo+9ySH+tZnVEkwqXi00H9Iv0yL08zhvgYJi3gtyBOgK7DERHDvmFk5onK
iHl+Z9agmr/Cc6sY8iszKoCxkVSWSv5UewKHpzWdzCOwokpiDCVM2+Gh196UZGCWnd+lFw6dan9S
db5h6VmbihrApDbfIwyenHVzrJapG9UhxiHqOzKDrJaqB81DAJ8wGyVHz8RZoEJIC204Rh4MjVfT
e9p60RWJ6eU4+URGVzGC2eLgLNTkU/NhXcZndCr1ULGLUG5tcxX3RXHxv6JQ9OnQbn7nFc37vLep
QuDJYZc0fkRH5JXCi477sBfwtU5JFZ0wMJlIIggMLwyAGxPZnQFpjKtvWoKB0hp6BpgTIB+8odYx
FgE7i2vfKgbr1OYFmbQBAPZbsnInrY5IOeb1Jq6gd6GylgsjEOZFX0UzcUc4ZPz1CSE4eWi/FB3H
W6Sbo+UsIyajAYk+KIe6KNERBcsy0jzogCV2TQZD+rcQUoOghV1FyjFLFWNam6ycvFiYXSvewKoW
gu+9SSIXRUa3jQVeiCW9MhpYK2Yss+qdViZ5q/JrPQDykWBXyxdq+I82C4eeW9VVBFnljryoXFZj
dNVTAde10/0x/TmXR4FgdqvARZzr12QXKc89FospHmNbacXWEvfbDSCM2DiJuQ1Buabc3dKuYQpy
IkmL8eiW5LtRD0+m9SZgVgmbO7jCdITzWPVAXnLwXhOEU1/5QQnUk9T49gginqrHeZf0HkLkWZ4x
ifOBXmXKjsl450ZTcF9vi3RTVNQ04/jNZ+6v36/SvGyh5bSegmceydtqYJllBezn0i/snFm2kEZf
YFyMZui5m4UytZq8lmlpcZzl51h7jY+rfS1zGl0Nx/Wq4Nc2NpkVZ+GLOSDmuvRH2dXmvUnYsv/f
p7wkjMwfY7eqexsmJW3hprFd6zVlmcwpdgsJvOvhj2sfK1+CSa9kZ4X/xawXcIR1jxRywLn7whRp
dqHpkYxhdYCnQdxX0uA96UjxwG0EgTwuPeIsTdE2zB6Y+lvi3VzrH7xXQlzT8nYHIGMwk7+uWk59
cGIkoPDm6RGOFxggL8AQeH1QXFCm1Bh00M+0t7wumMxD8boAJtXgpssGRDQXwCeTqxe3cOKhO4cJ
D4ZRkV5irIILHlQgQ8I9HmmGxmsjsk7Jf+Spa0rvKSw9cXjfwxS+3FkjCpA0cO0skkbR6nS8yYbF
7pCAx5aGr2KFAchP8lHBLbZISrfZ2qCrL7KiC2pxs3SUjQfkJkmI+5O3l42Fra+UbGCtwLuzZPs/
49zar1L3mct86ZAo6xeTkFF4l0U18MqlaIqO16jNTPxmbrp+xgfL3vBw072AxqKDS+6F26E7HtuY
xTYXZ3aX00hU8JttVI0JuZ15Q2ITHP/vY/5uaQvnv45sd3YZ7lVyMH9lHtdjwN3GsHWS90sSWicC
PzVKAIUxrGX3zWUa6sKrVzgWH/aSf+Fmvscgj/8hsmRRxGcI3NSBamTp742Terd9UjtorGJUZX9o
uUNshKuNx/MMbRBuiAWRUSnn33j2OL476F2yPwzAlijYmEPv57nCeQvLDtUIEmnbCQ/qOEvRzuSt
UNxTRjpXo4gr4napBlPaRK2G1QhlbPYEIJ96kCGbgOcvc/FlsCWZqxi2/eQgmRVd6KGIdlFMwYAX
bYcJmgTp15LGEJBazUEMEAyrLhCaRI0Io0tYuYZGRQz7BXrIdlB65SIL0MROZoEogn+nW1StefEO
v+fkKnc8nIYOfAaST93zuPHcx5+59Et5f9Z4n+iXUMKR3z9P22m/T4VObPosHU25OgesKpT0JhvZ
fAg3vy0UTPtmNvF6MIUt8P6Z12BNC+76GhDKQCexKd7UasUz5GAoPu331JxBbAECfa1lQvy355Uf
FwyosLZQMtxQsIoEDGdiZb4NV/0U5X1iYsyVRdwGDV91SiAlPfXlWbRc+spJ0oo4JNHWDGKJGJbw
jKrbnYi+fLKeYhptn1aESTpHKunMNwYIWK+ZdNiHnfnAVjgO/z64fHACA2tRUFKJg8d+b71JUeHl
iAYj3IOr5rWulT7mF/7MPgofi6fp6alDEtv9jlCPOZ2va3Jw2mdhcONmFLhZgtzKepWr5SIvIBX1
YAjYGGUkcCilugTd1BIEr47X+Q++HqE0RIHyuo9uuG9+sWq9A7INCozsjxx49R2Cemrwf4xgKZt6
/Be5fVTU9FEat6TZvnjqTq3zKR8LHVfvsUsK68YB6CQBd5ewhMBJQluv+JtFALTpJsesjCnKKEEu
5I48tWp5e+0A7EAXFnlDCKJkhcL/Dl3ih1KS7tlpM+wuZci1+iYffAggaXsyXX7obDR8TUMIbNU7
ywomURSVQHv+7jT1lBuFnwkEsAnNbEEuf2IdXnrkSImzd3teaiCCbbS70WR0zrzhRtXqKZQddhzV
lXXj97DiP/yWCPQjGjKATiN1OqoOSBZwATtlQ4iE/2MHUmwisz/POQchWz+wtHxMEMItx3IrUB6z
Jzq6gZI1tLk49twQKb4qbpq7Bp24t/pdqwliC33mRwjAngOyN9M1vtLlmtoispxHmIjQG5QTbt7p
zpdQdljvivjVlqKSfv4FsVY+a/P7TfSkfrzRKX09nrX0DRm83RtKfAVl5LMxHbDZBYuwbsE7hmGi
BVg3+XZfG2Dnl//5274jExlNwMdzbNVNoT1r8HY2+9J4s2mz74dPDVwTdEvg388SO1oJDryunbcN
YG6YgxQP9WvMmVPFzDRoFAC8Z90NJBvp/M+d37eKVfWE5jgmdN19kiSbBNXO5OTboxiaUYjZwF7r
iarxOEd1JNKZbAtezv4pfqjTXcfa3GOGzylLrJHyCDE01hEDGdH90AFQrxpzCVv8KEaNDtBfzsu+
gbYUEa9BHt8K5BIZ/zUaOkAOEcVfW+kLGYcI5co7Ktw3zX9xKhkElVOrih4P1ZTTUXGCN7AuGMXU
yKBNUmIGNha0Qbycrebt++IKpkm+MyWdHrIIsK31lRIPIWQX2QEcszJxLQT2e39HmmaaOZdO/4RU
MkixVXqtkpT5njftyGQQAt1JFC0b+k8nT3o1EHSpXMs7oTWevjPJwbdxOLZ6E+ASPw+C37IEdbVA
QC61la07RuNSl8qwuCU+NUc1owwQVjzVDbq82536vXrfRiL4gsYZjOPpkvhJ4KuBipPO8FXPtzJq
xcy17PvnTkCbX68ZD/BneQneHpgQDXXQf7eRDWVcWK9ZgbIvHfJe7ElASre30Nr86sVKGlvXUFKB
pIEAG4Y/pe8g9wSFoy+rXQWCRqifbpvv5HTA3zw37CVXsNZSNFxG64F2zqKFcniMkvXafyJNEI7t
AxvKk58ZAVfYkXmXrT0C8A3mi+XPBw3l+Gqiu6Hy0h1rFflnY7O8m+wqtuXm2EaMF5xIm79Tj8mV
GBUFJ0UOzt3Dwt6/4N9bzvSk0uzF4+If/X6d29VGVaOJZWD3n9y/GD2dDk15mdpuHrUXGPjyzIyq
gGFduNnasYptxLJlRat1LITWwxsTK/HFkV4/DP4HXGZG0FvGEeVAczzoA5WOfjook64j6kXjOYQI
wLs1k//gwVKdw5JssQpVTZbJwbKiNojFhehWXUhduP8y9zt+J1KWPqcJA9Qesynf2EoAaejwfy3o
P5wAbL66RPNtvGxuhAkGNZ1pAwj9aJxxY7E16udtQJVkEeDn1JD7w3u+jpEUVtaXFOgb6RV8h0lP
hCYLLDUDQCGjxjB2QxflGab5RHRNgpprlUdT/qZUKOOrmv0KsxUKevdoUCLfSFtHWQ658+rvEdaQ
u8D2iuZPZ9Ty3+BTJvJkb0CRwT0BCThz4ScC6BOQVCj78ATh3DHQCSc84cQbsC6vkq/RnSBdjbSf
rky9YlI4UudGRUorEIkeO7UszaPNv9X+pZTeU+Cqpye3yaZ5OtaNcKuYma00q1nDFIRslijoD8l1
KDmMaNoX6UEqmkkLaInYdACbGWYHjGFQFdzu+C7Tou0oUazoglBzTMtLWh7V4suMAF+J/1GvACcC
sRR/WywYwvSobRbWMvhxGiwh8EsWlXkbToXPu48kS/zNg/pcHPAixwQF2oHDXFpprOlWYVn6YlV9
cp+V+fNrkxKMIGqxirrJnCAd+kUv/LJlqBfcDxvbTr7wLfyLkHf8nlnWaOZgi4hWkqE931TU6VYV
U2C1Qp13PXuei3rFCeqlUW+fMFhSn4XlHBuBYw/cL7L9I1HjEUctenRfOQVancr1DdTc+/72LQLx
5JrKdz8naHj6/Hqc+k6fVz3Fbo+FRobMKpNBgZs9nDTKMlWr7kpJWvod9B9LBNxUHJZ2+cCZ9k2U
56kYVTGfNhLky4UHAhtCA13Uxb4cM8iBdEG9cLjwzY1Uc5NRW6aZ0XA2Ve3mN+kvZX1lhHdZCBmk
crUX2JFuOrsXmNU+lNnq2p2ZsZBc5/QvtV01Lt+Q27EoLDecWScYnm7wke5NtgOmtIebBtulkZWi
q2nsi0nzQ85Qr709OovOcH9Bw+ubCae90hjLmuZAk4DDHf3c8Lc0LNMUrKIvjkqA5yQ4+E13LgKp
/sTX7UgWShnePkIZ0dMli/67/QLlPVi/I/UkrVIbNWGaVYXImjjOKkjhAUlI8SZKr1ZzsnkW5ZWn
HH9e7pmVPl8kSn7XLO3aIETHVhyqpNmz5UpXBJfJqGJqfF1UdLii6McxJEa6zinc+B86+4QrOFv8
Qm/8YRPTclAPk57rx9ACkk4YWS9VdFAFJ4E89H5IBm09RCb5QFvkH4IUYdp0b3uKiyROg0OXiAJL
UzRoYGM8AmqcNJSeOX4jOtca5/Dt/QAAfE6G4grXPAnRN8kOGVft7t/qtq/vwUv7qlxethNtocda
Wsi0XVU94tW5qs6FxWTyy51aTPPY13tlXzY4SDDV8ux7yXJgDVEqoENXIqHu+yHZsgZpRFa1yRc0
wjRhbVW1Ky4diowAXXK7KZnigOWSWR+NsVejJWc6NtgizWkyO0K/MwI6a1Gmn6ej8UkCHs24adds
mAF7eHK/yJLbK9w01mo7NZdepQV4NnYX7upuBN6COvm+qzRvbnvrUp7AIGqVMqUCo4w3mFyBTdA+
VRBT9+WHXwTjFJsLyIRHHNE5Kup7hFrh9rZE5wQ4ZfRc3+tZsTy0O5mcB1FNrtNBlxqlJnD/xwi3
5R/tLYtyiJb3IO3BZzoHvKumGasPb391lISgGyPQFK9HbmCDo+sv0+uPIWym9R0ReaeI+og+Hvzb
IzzReWLBmPkdUQHisRuE6zQepaegSVWITeqLjfoxlKBcjAxjrVuI7lVNvoxUgROZssNZAnlpI4t9
0NiHxFC0D1QboD0Wk1gF3ibY7cjeNrS5FgDYQxctwtuqg3zOOEmpJIVq8xyRkQn8RpHU5uoXzEGn
XSQQnWkvb+FWyQgHytKbkiGpE2WGJChBcr/zPJE20vUkFwa6ZVL3RMTuuNwBE7SA5i36XNAkXpl5
w+aGbsbPGuJIsxQtftIMR3ABBCZqaRkZ/OlZCXBcxmv07IUYNhoAkBOK0KzxMHyV5Z6KGCbC0gPc
cd7WTSVgacoS5EfqYpH/3c0RZ2qp/calfhKKtWliIt4OlcDGtUG1Uh+eRC6lKgwAuBI7b0jvZ8F8
rLWVS7FL1iDD7HQRQIi123aurgCik6eFyTspltaJ67f77FD7SoqyetC2e6962vlFIIt/YmYjgIk2
oMe3fzLm+UZVY8p7EQ/WaqRvjQwQ1rHl9/7LHIEmjvXcU0G6ITAPSIa4BwUy/oTXVNwR2j7l7jL2
6BLDm3GV6lLaGFf5J05kg5HtSFrbaOk+ijg0NLgVRH2aNoIiFywCqDwLVGW1Jrbl9VCLTmvmfKTZ
fuiRMcLPpuOF4JDbKiO9xLObIC9VFNNxPiDz+foto9oxa1GScJTMD+63GKwanpk3HiDEK4myCKa5
Ed8TzzsR1PS2GW6ALeMiMjpapPv23Zlt/ruuLJaZ682QbbKGpBPZabZ9dlQVdLfDogTppZn3GRru
yYuWuobhirP+1QJacji9tCMCtTUXUd7DA9H7hZhMUmRYypB8B6r/TTD3z6mNI87Q/QpwOzFYVPeF
B0ITxgFoL/t7YgxoVy+oCsQBJUakBnfuNNbNj8GKdGQb9G6NKuK7NLTtQRYJfNcTIpjQUzW3vufa
1LbjIDZo9Onfw1Pb5HZ9iNJF763YUVEwxa/dMC6ntYPTdeibS265JyAhoTpQLSIbhlw6sqJk8F/8
kqEOvlr0V0CksM4QKZnMKn0VivJvjAJvzOEob77HicWtAzwT1a1htqTVbIaY5tmXJha2jTE43JKC
al7A0vIQ9SUgX7c+RFW1hQl4sa1YN8XLRVKgooBhsj+UbWCMnis6VWCpXZLFvlmJ0P0MzZiEZ2jp
mgRFy31QyimGyUs/gNUiQDYmHNFj+x1rWjVKSxfAC3+46uw4SPsARTLsbEyPiXu29fx8FaNFj2cg
tkLaGOjbjvAKQYa9fhJIWNLMfMOjyrXZ/RWXsLjw8SrLi6GqoFcno0aJw5VQeUYgy+CZVhnUmyAK
fsl2/MMava4FSC6FXgG5HHCPwSTUz5ICn4exYjrY/V3P1NX0UixcD9GcnVSc66kLfVT0wWzjt6EZ
xoAsRfgahsiQ4tou8vNttBsbJycLDjPBuWRvOsqymGl0KVqrZqXjvX1kpLRfboAEHOvyvIDSKCkI
88k75bri9fV2vOHGtpJwre35wCgdPzvfF0AMGlvBDV5aVB/mQYd97Bh4u0N0qJcwqCVSq1d4t94Q
65RMurdkQIeJh66CGxXuXDxH8cmqG2D6PVzxDqFjF41O4P8Fu1LVem23371uAehh2KE3bk8qe5jj
b6iaKDLnJgn435b2TSsvuKdV2fmknL3A1iTY+UB+UkIJie7hlNCjmZR1ULBQZVLmux/0F02COr27
bFC7USnR1hPTs66QUA9Go5hOpTHkloJmRQUXwwhEmfn6wfes+CflYx50hlz6RVngmWzgWthHYGPB
hiiSEQZJkJmcJUY25U/GRG6MISTWvyKMAyCBez0ZudGiFfrxgXmkLBHR1ptnMkIjne0tN4PfPif+
x2TORw/83KkLK+0cxck0hn585/OC8Tye2VPT35Zv0sg4pZgByP2P7AO0vONCJ9UV7SZRQjzjAJj+
fsf+8VLbb4lT+VKW2Zrtgx0JVJnB+rj3CyP/zPE/ttdOvEoOdwYn+3KVvSzAEWkpdWPp5BGJ/xTj
izPp8MMBPs7jjzwwEPwnsrs7ngk791De0NzOqLJhDEaSfNZSFAgZYsJB7dDMYEt1rZEVkIkNXfOp
ROoBPPSCQgOz6lOy/tujdeaOGXy14o6QOunj/kCvXzx3Ik6QPq9AiZqGvLA1qPX7n+di9D7THBBg
diFNQc+00BYaco5J+7pQ0mR7nAqZskkTOVVDnLNypE7BXffhsMnh6zdwrsGFKVSlHSQxOdTVC2ap
cotKozvQroeqMulrtm5PuSymSDmBp8lBj4ugJSnxw7tJml0TTnfZl9s9tg16LEQ/lh0bZlV8btnt
yq2mAMogFT/hVKJmhKbBYibOHryQEVY6ItmCHjJ97h1axyH6oYOT36JTu/ao5T8x6QPXEpTArKk4
+8WdGfbckdtDdhej70Wwsrtl/G08MXgxq4zsWCHnZdpiafJ6CONl91hGFHmuDwFHGxZHPlfsN0d+
h4c8vkLSqP9atrRG7UWcDv7KFmAPt5Lll2y35/UTvbdHxrIZm6Rq99XGpV79dCk97VU7CvwyyqjW
ftzysYs8wY4C2mtM+y6fJePhjNFmwgVGhX6c1CVeDsx2PfwbeFC3tuH4rMShpmU/55EB8uBcUBnv
mYD9BW261gh6qnX0ootCxzINw8J3pYGBNRp8usdk4KqWFpIz8nIfVJ7d7Si/YnT8d/eqRDoa7znj
FapBgSzxk46OemmarrLiGLX4eiewFkUGjyB3zkLGH8VKshhSnFb1WVido2FEC9xnppmySNYAEiHA
9R6hx//wtrufgHNyVM8Yv+7thOsUNwiozZWANnU0XL2TR8hzM59eN2F4AfxbmS9hBTGGw5t5g+r5
2rRo2DdQhwu1GMfv3VfbFwShP3GXMXHzTllqBMaCSHN5u/av9biiDNcnDQrnilx0ZICKyFpr0QaI
TagxERdxbptL14YBZ5iDgk/ttqykb8+zaG4309q1jIxyY0ko+nNIsP4mxG20DSi6ofPl5ltawnDz
w+ukrhXWis9PnQKhsDOjbr91yXLfqBnKJ+mDOy/YHPZK5mLhyCUudXysa/VKdgi9la0UBM+Q03bN
qoSKJ/3vGoRgvC3MiKdwveETSmoT3erTCjZMDer6w5c3aIG3z25FdWonORSI68LldXsTmHeJwx+A
7TNmWLyLXSfmE6lCdCA5IZSMqPvodzUeJ+lF5ZmrIg7IM0dlHQLbVkwuCVjwklaGHptPODBJKa5P
VMkZ7eZRHNQvCFIQSH7PfUV6/tkfEOFNT9AGUpyylWxDPlXarWIq7EFdUCsqbuUX4aO3ivXLcdBo
8i2NQ1HH1CaNz6mRfcFBiqiWCOHpXtsH53tX4eNHrngN3lOsYe0LDf6u9wneMu2Kpd9u87n3x8f3
IqDlHRMxsmFPFf5sT0LUSjfNQkKtJ2n6xvbKxNxpvZAKIi1NN3ht++joTB6HUprnEdWOFoFbNE5P
YHhJ3UnIjhqtsFWk9YsMbyso/XBXXQKn7USUdcJXcoDCbBQHEkU0raczq8z87vJv06neHGgRZy+H
5kY7vqOW/2sd0OeXWWg7xfp23WXzgNE/xzyMOSJMFuIeUXOB9CsSxdvq1JmAHXCzOQoSBYXskSFg
sZQPjv+5ZZB+tZCOjd4MCBTWq82STm1nPeKr4T9d2s06Sun8FkCgRbl4NCxvF6f8EM4qj1CK47O9
o5s234GtYk9Ttqc5gKAu6UpkdVf18/UU3cTS9RMgcL76VlRTCS2fpOjn75jKQyhQoiR3osD6aaY+
QXRtfvVmLzhi+/5ArKkk8VsGpFVZyC6EA8hIjJK1haD82uj1VQjsmQO3d632I4PYZq4JFrIf5THQ
LQe/OtnVfYb8BZIPWOwOHNw289B3F73E9qxERDy6KVdG9NA5VIhlRILvrhHYOmezOHZtIjzKjm4c
xs2aTxjJTKrz1HXGyVGkwpCUm2eWqBzeteTOPLHPJsJeH0xLdx/gagnAv3jRwzOtyep9UwAjY0pm
KkVXqPdgvexo3ly5ksarLZkOULHJRusdWQivefDV4C59B9fKYSL+Z/DVy0HTZq7OhGEwmEl5buZ6
MEkvroE+ZreqODR1OXDrh2AYlxytcjTK+L+NkcZyMDSuQ98iYRyK5Ny14gEbDEh9qMRVigsHufPU
+VK/NHxaorpmKGDXM7J9ZZI2ul07gGGhUiA09sEy05tlGYbmchjjILPabt3gcI178SnEyB0ErCzW
Tn3z5eEUIcuKgVjb2/oMwBnmpxeLxOrO7apHULwWfD9GU4/wuwbTgIMGrrfkJqd/0vOTK9uvtPGi
9559fBXOsml41rTgy1kjRGxOTzxt9ModG0pWfTSzMl0SJPMMx+4WO7qUX0EkQcMruD0kA1bv0msa
JAlA+gHeqdEp+0sWUHIw/ez1/kEd+WC+JDKDOPfRkM+kQ/o96n6QSHfkr2MHe2n8xmEIciYUOqvJ
/keiC16PjoM453L8HgHWqDEXtE3i8ezkrvzJvQHJK2aWSyPbrss10BqL5akWnMlZBdYxxFjpnfsC
EAkcmQb5B5SJ8pyJSnp214NnH5LtjXC6Z7VP86J3svEr4w0p/T2p2V4cEi1as17sxaGMx+mIPSZ6
MBZGLoQo4y4g8UCIURzJIBVasfb0FFWrhLJEbcu8Fc1gDkXhwxnM27JkpLb/P371AlBY2KAboMO5
BbCl0mPoe9l+QU8PY/g7z3kMkF82Pke6VUMHSx7ml19Lix4HzyGS5Wxd13x+kdr/VJKi8fgR67b7
59INgXz5wn6kMflxjWUcTvCXHIAZ5NynxZpPvCxqNroIdb+tUmmk/AAPR8HMkI/dFKXF8rhyOhGE
l1YmG5Yese8fyU1Oq9o94dS97ijHUFzWRVZHxLTcgcBsYZzXQ0BcfeszJBH3zpdE+zicrlOEcNj7
hIkbGtlInFLn5y7zSYY6AMFjsgKg6xBBqRe9m+6ZTb7EZS3imunvzT3NqvzSxIhnq96pqqEI6yRR
l8CZBbfh6Uq8EjO9lX6Jh4v35SXDH6RgngDh4yH7CVcxzvEmazelB5SdyiwHqrbYgzEqQ5dVuYWK
F7YXi8paNEyKML93GWOMDHezi6g0mN64gyYe1YGJ73b2C3O223iaEx0U63uUjxXvdDHd5K2zgm8L
BXH41Wj0jAtxwsZo2slr+xQYzi7rJ4F0DzjFghNL8bXRqWBby6NtBn15ys4sBipuNBX012S2Yv9b
j67CJ+AfZXP6u6Nrm9npEH1i31LPnvDdkbKJOjSZXPCii2fdAfgLfEllM5yT4SCjyPR4q8MjAhQ8
x7eatwArgJXhF0nOaT2Dyxb9Tfm3DB3gBXKn5Yi84o7tibzbFDC+AkhuRVdczlMiqUKBl9BVLeDj
LvZJWTszQ4F1eX8xK2E5/dNegCzM3iBk4+kM6dUKha/KHHA04jGU5/kCwclzRIPNi+YeQ8X0px3u
wr6xBwlW7j4M3zLdzLXxS/NENesBn/jhYFXeztOhguMtuTjTURvQsVsvZ8RGy/JaUtMvnoD9vdwz
MRzpN7sqlRdYPLYfZLSwkNFEiekhGDFLX6resYEjobI++t2LnBLR3XyQs3z8NDiAhQzaJitzZSGd
9ZUqb/TnUxVO1tYy6kWMkeZpW/IgHp12OoY/Cho2B48QXa8GxtU9iNC4AVX02NxH5dXDuD+HO8NU
K1IYhDoM9EVx9tWaInV9D+MpuBfe5MaP+Zz1OnYp7gfCBbQ0cSC4CUxUiIBeSL1NnIeMBKJUoNfs
B6MnJAar6bqJ4h+hT/WJKrefEJh4saX+7BPyYb77tBmt0mVnxFmeQU0jTqCuqep/pxK96cTEMbAx
x9JgooIfxuQ0uLGAEULOq1OCQGPi09nZWbjpqJ+wowF0z6G+5uf40OUHLigakhtgFm3O/Bup5jbe
IbtOw/nV7i73ZH0l7Zmst66C5Xf4XWOht1FFE4bfjafs6Rays3gN2nerOybM1yFHyyhFjhzAFBNY
mMbcQljt/sWNz4OSD0peLblM18WOnRpjdiHtmkSFVbfmGkM6zAqyCS/muNo8c6wa/T7nUuv9xw/F
IbI7DZnsgFoaNFSl0G81xadoFsH6ouA8mW/HcNxQrUGdUGMCRraXzn19W+32mfio93OSRspqCci6
4XoGEd9scQKH2hM114TmlxFedqm+yJ34HZ+ZPLag/iM9LofOjrzikHMOdmZP68vwF0vD+i3AGNmz
SKXBT+HQzDf+PiyglzdT5GSFzW8dEy0zi8wKEt+ukD203+YqoDKpkDY2bmU1vyaIexhf2738nCWD
LtLXgZYff9UQx2HOdjTDi6aC7N8PNcJva1jlzykSp5uAFW6MJSnEZkGw4aDIz96I9QnCuZl0Lzr2
Tg1oGyqJJQ7QB07IjWM1cxQwy+7R0CUkzxciinRm4j8imW7/xxBoh+zSTqhkAWU7d0P0Izj2lSos
6GmsfUsgjt+q9NByKevyny0Ny6j/GuybGsTvhlIUi4WGxoQ6JvI7k4mNRKC3o1Bi9bGSFIBlsN+t
XOAszd2bMyysS6FniDdxTnb0gvV+UUNPgIfC7Un1pb2zxojQdPH4wnxsXuT92lNgeHcuz1xCUT4e
wsnxDfQKkDxAnI8WJx6O3PHm5vOI+Ft5sMHE2mywhMTwUL3f6WJTpzQCzPYkZVn7mZxHsHS0G8wH
a+ReA7NfOM4CDNkfK0cuHDu06TpEuaqbgpU8WxvZ8/zFq7sCN1ZnbmFrtKTUGAs1VK62JLmtCmUr
IjI76RcGrt3GZH/nZKDo0p2H1MXkZI6gIjMYz274QSpXdMpnWCF+F9k4+mijjPfzN/WQkWe83GWx
ebHvzgCP2PybEmUEkX0kL4oXYZAI5P+D9WIbCSwdEE9YS+v7zvZqHkjXo1QI2K5CYY7GtpX7Cv78
lkaaUw3pbmghGkE+ijMj7AVuvUMWk+Hzjr9fJondq2747oMaAOc5lVz6tVJJcE+i39CJZaYcwyBe
BsdNIcrjTTVS1NV7atnnp6SSLGCV8gicm3ci8tX9mAtjWE0XF3NrD1Xpd34kGtbfbsyluJvkFFph
rBMjbZWRbSLXZyGOdZ88NXCZMwjYm3zzqKS9Rvz5+BmhZ7KsWg2dPhFIxcJIq3Jym8ajyabWuinJ
9L0lNomkZADNcwkqTDahBFDTXxRznxRSho06en+eRC8luNBowqKbEjQLdETem86Jv5SbVZspRTUm
i0mrr/TBsbzdpFgt7SqMtgQi1mSZ72am1PfAbicAmvWNpd+QpAeqLCYmVdTFPXjvytCgHmPFXpw/
6j9DH3fzX/zopti8uCLaRvfMIHpup50BTOK0tFORS22v4IifFfvtWQwhiehC3R13NmSJax60YB7P
/5oH+NKIZK+Hj17DpU1vo+sQDGYLRNImp2BVou2tKFtwzZIGo9ELqfBKdzvj70Mcmt6nF/wOmtcG
zmTO8dN1yBumQoOEkgFRmZ4wfZR//cnVEjm9VktOVbPvECAoAniyN6FU2kap3N+7aCXrPG7qLuGm
qm4YKW+owTItYhCTvFN3Z2XcmIX6wotNbHkdRduYay603RWfD8+/VIhcPVA0qMLgIthMbzg+h+Sz
q3apS+ELZVomD2f0cAPUUoQ6+2/vKq6xb25cipeAZAWp7mva/jFF9HlocJ8J32Db0Y6Y/ipwClHu
nYI/UqifPWE+doQKdWI2SgFZEqZxfDRFr2WiGy3v4dmI/AMfoVmzZGiAVn6UL4JDl336vMFgXlku
sZuvubELmSKs9kfr+MhsDkvK+dTS1Kyc0KSHD9/6FAKoONFY9wyIKHTcA2FE/0hKXhSOm91DCBih
KAt3n8GkXmlacjo5nWCDHugMelXDlgOki2Ze4D5Sz47l5iQSpn8Gbsl0EIz31nPL2yH6YMO3V8Ox
rAl5wnszcuIZozAFF3Ygud7C9XCpxZAtmU2Wrxs3pBTe2fXlLixTSE2kD7mCyoCvAQorygrZGdUi
oVTt5PL3UMIBcCSPKbNjQ/b1jpy9rGyTMg2xGNS9mCfSdJP34ZM5B7UWBO3z3CScNRhYdbTYa3LI
qcY7UVcUkw4kw58xbEitGtFsmJ4gc+74S2vPe3hQDhKfe0y9TLXr7tZ7RLdbgv/JwSuWOp+l3BJD
Q8M2s6cmMNks2GxoVTYjO2LkHzaPfxwhUG0x69MxQhJed1RZPNszOzopCV7wYDnsLxY+SpKAaLrs
juBil7n8pIlc0o5ZZO5Hh6/uyy2q1XGcNJogVNDUN2Ts+Y1pv7TDipuhYycdWDtcCqpp6kNRxk61
TS62NiqNe0zwsoZ1VW1BQrau6AYhwf+HfblEhZtVpIRqThyPcfWVoxOb7YznEiv1YpK62VgqWoxG
N0a8i+rpHN412otIVEvGZd/saCk9iJ4nteFQQ8wTVlszAeCnXZw8msaSCDJEywYKhYWoz/qh4jeb
+FlzIKTwAhVetP150i4B0siYlklYldtojexNDrZ7Kukx5ZLvllDwTtYyMI70slqdoJOf/9v+oJUw
cD17OpB7JbarF4JlrA9H1DIPXYnCoJwY7rQxj6XwRNMOel5sPIiOYdZi1LyaXexX+F3+pH69m9aC
Fs+tGfWJG5Pg5qEs65i0ukz2Y0bseJKrX+S19TWEn4IJkmudj77YWYaaSXuO0rrcjCT0UDKTFKye
NIO9XY0WZLy/M0rLUli1pdOENUocoVO6nnkbuVjg4c1wwTmR9M1CqY4dvWEZ7bIaK25qxcrwOPFF
/cO1c3nIDhvIFzuNo/rKoU+i2O/wlesOa8EQfeIjDWW/ID9ywzgB1olvqoBrYoy3k3u4kDPIOxcX
2I8iXI0+7bwxIHab6+RIEM8dfFtUrQeTFBXuiDYnOY7vHVZjfRO3YpEEzxrwVS5iMx+zKKgLUApx
IJoTx8KOzO3hr8BrBy9RopATESdSi4pQeLm6THj/0d9yqfcB5MWGSPYvEkP1qJ/44BBczMwb7/FO
B0nPJFP9VkiAUxwutCLhn+vGCgTJCNRDaBQ46MkiXji9pvbBtqxo9Va3DGjg4RYuzNRkb2CohNFq
qXZrj803yw4Ezem0jyp6ChvAlLpBcHBXvSjVU2GZm7JeyWm5xSEJQrdRZy3qjIY3Y6dnmZv4/QWi
YSkL9Kz+Dvqqd2OUd8IosvVeX/+kbTr9pr9CHOY3IB/ZGYakF0CXVVIKeLhslSFKxy65/1OVxzsL
GNAFVCNQpV6+wfhKxJIT9D/KThDezmtGGFo2QO9vrj+69NyzT+8AymUC/TAgw/Urwh3sw+bgrNR7
sxd+9LKxyFtNM83uEHZZjkT5uXVal1XiM78SOGa4nHrOsINVlDkENf1yMgRnSmtGtnvUMUIKBzKN
QiFTC/SmUm6b0Ge+rr1KZGVo7b8KNHXLbTyb52+8tOAhjb5H+gJNQkIXiNiyMf3ky2DKM7dkAy0K
gLiHNuXLZLpa8HAzffY7yuipZZW2ukHmMQCPTEz0VRXhzAP4k1I5kxr4rBdwmIEA/fzq4D3/t2fH
wnrIfnfh1W9AqC96FPIXNk9uOHo/ERqWsVHy+mWdseQ+xGK/VYjqmgN2zYlX1HA4D4U5uXB44lXE
vNtUoU5rnzc1LsF+YVQWTTGCHc6X3Voyogt5e8hEK+SDeuo8ql5IaNT1V2xTF0Z+Oqk9/TV1Hxm9
sqFwZpPSCRYQnL20X1lWJqqm4FvotK2hgCMMdZ8RBYS+hDyM0ZKcwBNYS7s/R0uVbm+2KVFeFSUX
oFwhv4GaL+BsJvtTh14pewrAvimLFVwwvGFD4WGZ2ZTgHx4WYkzKtKWIBBrX3AZWoD686fgis4m8
+FRJSl7CBnGYjgtVh+WptEJePNrV90mK44Oi+PJepfuUrLWSQ9Bou8DfW1tBpvJVz6CMANwBNWN4
UKST3k6mq5UiqHE0sfcVJ34zh+GsCzj8MsHBaeaceq1OhPU3nskARv0x95MXs5XwKAdhBYxSfIsf
tu6Ry2nDNaACehsu5s8Fwxo/Zl03b11x9ozNNKyEkD355rpdtP6IdZRGFIDI+44WVPabstwf9MdD
7Z7oE1IUSn8Ecu9bP90Jv46ikhIX4+BTo/uT/tsg9dENdkGZUugYeaoC6mRtZPkgMwyyDA/n2iRc
IwrsuJe5HQG5ubm/lOS9pPFfm9MBx+SVdsyQxFWuTKixZUrQblTZeFe219t74uUNB0UINiZuBJBp
JmiAjKJnsfR4RrkyKCy8dJWMKZs+fwZCkGycaxzAK6drjAkOP4pBAmPJRIbpXrp7CzMMmvBvNogR
/HAST+BiTDvvOlTf+qJ5499/v9o75/pNtF4LqbbAMtlWj5KK5+adziSuDFxDqC54cxyJjtNUJYYY
/4G65TTH82QaaIaYJSv5bCz1hqB2d7IXPqzZejfjjKM/kBvG8pMACZ/nCAhisGiDzIkbi0Dq8dw0
GjuuK0fKWc3xa6fUnlgpq+xpdJ8Y4AT7VmMOqAZ//zPmWtVvQxudBY9/Jg/l3kKtW4C5aPkszYG6
uc2WuEeVTslESXXzrPJYTnDsAzttUD/RvqTGw/lCrbW8kH8C3ISLAamC8/+0mxKcuDUxL3Mg03Vn
asSyplbsB3Fer3x1QCP8szbMNFqPpkERM2fjdz9xoUepiGSf9+VHZ8A9HiNZ2WkMDplA0gRsbbqL
5YdIaih6fTJGF27NHEOjd4c0FMtZYA0Cu9M+IybNh9sH0eQAUnqEQDJEgMFEysHvk2Oo+LO691v9
fcOsyev8P5U00KvaoIiHztPRvItV5eccU49ZfleDUPmIjQ2pp/CydnnplIkDaz8ANEG/Lh7GdSsh
BYBLDjNqNZIUgBqA3i/Qg8oVoWSVXRFaZ+0nYo45/4+O8K7DGdw9p8fRBsO87BbXuc6rjDlA4o3/
3iI96/ddML72SSKqsL77N7W65TXSJxnUkeTzvU8YA7He3rEIuV4vX8179th6sN7ejrQ/O5k2hdVP
JJXMQwk7qDVn1eFeLk6A71jYd21Z407hlv0LGkkMkR14790DjSN88yWSbtO21O1+lB3Xgsp7SZRo
JlSZih31Rh6Zbm0mCviWjnT99vk9iTh/UyS3CXn290L6Tzfp0/I8Frw0B5C02AjDN2/SeSE/OYAl
mfnrXYy9eNbdxNuqrU4sR+M4FoUPnu4KN4HRJLbjWI99yE6C3s9C3r3XvFtWVeSGeMJ53IbRg2RN
mudc1U4hByRYjBM5ddez63i1S0WG59KkiK3z1//unpbHsvUNwu0U1f3MRAVa+KsJQGkbOFaxiD+R
Z8nzsqoA+6knEhpCmq/yHJnpwQxQzusmt9vzZPvH5s45m+WumUIVWWWG6N7Z7II6Gn4geIDPMf6q
dbyga2BH0VkcWIHslBOMcwGuZGS7HJkcpnDVnJGPAD5fpxmNIBkHGjXLiHmBB7CZGWuzWPuwem1r
a5frQvVB1TYX8Cq1XN3Imxn94pBvvp50F1A0QRN7THYiZoXnZQaR2lb5UVn7E1GkAd3yzSN88H6n
ZlAvUCOFMUFreEu6Fpvx5jNKvqY4VVfxySxdC84pYXVf+VOLAOoL2AGT1tX8Sy9kuh71i8qKeVKO
Jp02oAKSupK7vejJxFuLVtSmrSz2+bAXkDWtcvoNZnZHVrOA1xR+vKFyEKw5KnpjwbO87ygJmvYw
Kln/MzUMVoaDrwJk2xwg0uv6ZNp+YUkQbCmBwthUyOd9gQTldH7BC3OZMWnqyb9WPNMq7t7eOqUQ
q6IL828aUP3NzAIvX08VE8pzjPp1wjCkcNpJ4Y1eimFWJB3X+NoRVHNE3BWAL6XtpE+sLvG4CR9a
tsaovxw/dH+RDjLcHfez/QC1BLdZ6+qQJvV4IDaZWcOt4Yi23AuKLU0kmcygQZ8MNHRhHO/8ownW
oBJeNmonAuc5jjIRlAAZByPQTBevToFv3EEqHl1Fv6u42GGJKjpAgIsPdlaFU4aFc9hkKdokszbR
0P1D1uzVTZqKa1zkO1ae2rr6DDZc8qv8yhjniG0Xls8SAzukt6X8xhReerE5E7nRjl1hpK9D2QJ6
qWlceEBmAEWxettYjHp6kxeHKmbHsuPndDsABlz5ukbiC63F5uFgNT32XT62aAC8xiOm3Qj6r0a8
z9uncKwfP4LCncWsTIwVbEg+Pk45TAvauFxsQE0ud0o062ugz03t8dTL21QmIqzmYsqXWyR32+CV
qyW0gZjiRFameUqwziO4aIHBHCX3cJx6sn8w7qcTA4TpY6H7Xi+egiTPz+r4N9r8G9gqJTTYqKub
kL4hyKGWOLeZ99Zv44x/9BKOMMyoR34it/tOmt6DHqwE6FXy5/3xpNmJOfYZyFBDidowtlbziTfK
Dv4lKieGLX2V7zKQo8NrjKg/kQHSLerM86n/RPYA6XjcPgGtbjKSGgx7y3i4XGebVsOgw3v6kgQm
MjFYVGKaPTYDS5YE+zU/kJfYg0srERTiBeSvuUjAzPOwwBaivRhM6FV3wqs1HRePZOch/vcknP7h
ljdwenM4mEDHGFGQlilxPCYf/MxLrmGDe+f2NcedSWdzdUokCKlwV/K9WY9u6KaHw9Pnz+Nb9vsg
9lAZU4NAaz1gAkmkJVLtU1kXE5ZWF8fPNR3ctKGyMxOUMTwvt01a+WRnPJ6F+nhB8Lui+Nanh7nD
uepdPX3hilX0OQs3zCiPtvU9ZrUWBHAVA8F06Lsn0FhC3WrzRMTsj6Sv2HzbafNY5WJozzDAM2/U
83w9vBXISusP3qnsamH3s+1NlBucurE+rVg6OXFQ3kGVjXvo3QLtWRjN0m6IT3YJYgQKgBVEdUSL
mVmtbBCL9n4R5sxi2vIOkRYieIcxgOaJmZ9dh/++yHwYjXFH/FV8nN/2T/0X3JYhM3LZCTrnhC2R
Dq86LLmUKEYFULzLl2Pmx0lmb6nHuREaSETWmwHKdkiHLjO4IK/v2FUeioPY/Hlzz39PIt+8bXsm
KUwHMt5T1bLgtuy2DrQVk6vSONvNKwG50ITSPuNCS/6IkXz0kuWkjwQ+Hbtjo592cRcwuuHu3DJW
QOBB5gSOUHOB/mKjc5aJzrpOxzoQ5x3+L5frh1w2HMhsKyHhkLIWHwmQoPXbaedFCN2rq1bszh2e
lfP1paUQF4XbfwgjtD04SMNb6d18GvBixX9p1sYd4vLCZaKsw33nYsLRHNICODp1xkW48d+2goGV
QxL3PlHp5Y5docyKDGzrg5Be85pj06CZ0no2C+aG/lYCamT6fOroPsS3+TRepGEEuY71p3tzJ2Pj
FTQVN0sLLAL8vB8mPMq17lBuF+K5/W0HnLx3jhyfygpeRamLOO08sqgAzXnr8V8rMjZ13CqHY0vl
+1+Zc8A+C3nILK2EwrdtncHka/zNNWutSNQzKakjsQnMNsN8gxpzKDwPQHmuPiq/DRT5HTDOeunp
koyfi/hdO4m5eeyFFyAkKRkIptQ0TMIirYP4ndxzUlB4C7gUuYCFgpupx2ET+dJJH1OJosdsd4yI
aM8EQKmPQj8oQ/sh60//O4aSx4Hxa694PvNptAXcOOFr1gfpnlsoyYunlLw88754qm4rrWBPes40
ct8+jqRheb6RIYFZU7VRgae+HlUAVRHjosL0tpDLbw2N72Ve/QghIna6t1y1n8DkwMBgNjw5blNS
Asv7NZ9S5uey2GCbmrqG2O2vwzBVqyfarcf9kJsQdKX3zQGC5nJGlkuhjdEUwoRBk/rK49prb7KL
la0CGdTEik30+0SYBuYFmII3XWNQ6zjb/af57+mOxKww6e+Wh3TACQF3n94wF89HdQN+oCzAD5fL
H/YCBAfVfsTIe6yP50FPFK0EkoEHAN9/Ssiup6i9/WuYgjKB9FSMukWJK0MmJCBqtRkMgeil5A4Q
jT/+iIUAiNZVmMUOue8Hn9xCqnaGegTOv6UiB8bbyZY0i90hQRF+jYCDlagY6v2W/s1uDFkk2JlT
XblFyvHLaA7Q8d/uKU28jHOHdwYwkAI2fOLu5/3qFY/hJ1mfvAp/XYJJBqFs+4+lFS9skio5IaJ2
LfwnI7ftbm98BrTZ7fTvU+N7C5g6vARvNxp24qyE1URR3PNk1NLXj+5n/MA2OF4o+fB0dVmLWgb8
/Og7kh3afnFxy7u2vKKwBbOmAJI77i5HXSkGFO4CkZKcWZtzliqKY1O3v47U+nIxKdIaeL6TyGZw
/S7DA9o0h+TanHC7RHNF5sPUkNCHSys5M/Bj824yXf3d1EjYWXcuIxH2hu50h0mmSwyab3cZd/IX
hfNO1PQ8UWnb7fKQ8W5qtCNeRqsPhh1Z7jN5+ndxJEePv24kfozqkAQf6TgLA8m0oUJ+J5c7jIO+
dXcbOdesthNd7DQDKy9bMbLPZRukNs0lPZxLEVbLBKkCDRH1YHNswexAuhMdt9x8PVEWbGeu+WmC
fDb5rT1Wu2O4gLKQ3iA+CRiWL6SShN1Sm+CmIwpV0ZkDCB4pxceFpcZlII3nJUY7r1Yr12RwCUd/
jShHMP9kfjMnvfbJY38jAAAjYqyo3hAuDd6WrJp1jJk5VvFiWfVKge+TP9Qw9sFAL1frE56JH0m/
D12/PRLlXdWxfWip/cF3IT0N+ofZg0hM0C/eTBR/CYqa3jYhiOCWrJcY4Y6H4e8pbwWbZ2upCyGt
z0UcbPvZc5VcZiA/DMF0JS466RY7bpkLiaRORtGOIhyQIy1WawxUHaGW0gSlRwsPKcrCDPhED099
8ajV/jYcpABV7lDXJFW+iq8xY8mGocSnc7TL+VFetq11OPATLGU23NccfsaERYiBOjpRSfF+25WP
wISY7tdIF5NABd5XnuELF68Nck+PtmKSQns9iD5q1IGsiENOw+W8e2AYNBm8do2mDP+YK6SQgMBp
XeADQpHnbcly4/WEJNfVjW+0oT5TXHe56PP34i7DZge9G8K0rzQWy6ytRluqF0uE4BQ2gHIYqiS3
yQf5j2oUpjsLvYiVxzYIj6mjZDke5D+OM6qbnTWkWM7qKxgYQbOHOqhxoSddmLlWpmGZxy+33mYT
w1G+urE+TxvpEdo2O3n2qHKt5UkiddVXUl41y5AZC9sAjbaRFkRwn/p6msm0EpacMs4DGcwZVb5b
KUXS6xif1VN+dnM/02BWQ+j0gnkX4eprZErnSnl/+UusHFFvMBNwJx3OwzbnmJdAxfaggs682LxP
Hn57gSsVZnAC5fseeSgBqLEGLLT2AjhQ197N23qehBNZ6AoGT1JzUr5wJPMikIi3BTNDKAwvbgYe
kzfpYr3EfTUuvgWJlzaGZbTxGcSMlxJ89GtgxS6jZse58eCj2pNbRGbnb5cVmlFRdhJPn8erlrJb
5ZSrRbH2t9qLlNdNrRv/wHpP73Xz58MVnGSI8/vUsrRxPk08kHKAvkfHiNjSY12Zy+SPJttl1+gp
K56uQCCzRvOtqF681oWQwZusYUI4SQxiHm1ctsGR53BIrEtkSbCX2bgkW6egHwkHbGYSvC2seprg
6XSv1l1Cy5ocl81bjHSm62b59MMi1ZxCLYmhszdjH4dcWy2rLpCxVdnKBIGr0h8/ojPSuaeTMKKV
iG7tMkEyFcoRGJK9Uux6to6bPXaEtwdpwgWHuFovclny468CR9xLEKUTF3r8/zLjwd2TN06bnYKn
oDgJNIT81/ggmOvJpFJ37LJsyXp7MiUYrsGCBusR55s5zsioyxlbEXqn/0K3OCdrTnyUcSFsRlAq
D6XtGSsyDGElD512tkJm3OUTQDWqLEADUA0fg7hCsor78a0wSZdDbOUP7JT40f2HzY6zJQsClB1K
/xbOTMUQ3c/ff/nGXJZPyHIrYfbVL7OpMFIR3NOlmPMKPk0cUGUXxNPqRHGnV5iWlGKDAFrISzfU
LkdPmPsRXdHmk6Alcbku/9VnQcZwIw2jD5W1wdacxOSamhPEMKkwJBMtyIlODgIg5HBJDre+cRFY
EfGx4OB0bPpCNKl48OHBk5FnOmt6WdL+rNoi+NkwSWztvjKWSrIVvhiK6lgTO/85pPXvxkM1c4CX
H7HufFlFM91iMiCznilqTG60WK/9ms7i1RuCN+RzasCl6KFKgu9wot0841atzSJ2q/OYPKuAqCux
Ma6guCrJoG4mdDM8zstYmsWIzzOsFnu7K1WfXifdKbAzbu6CwHZSi49nbuxOWXXD1G9CwjepCzBg
evDyhya/TwxAVViAp1MOl57kKktqzICYAXhkc55tv3W1TjhN/oUtPNJ28kXtvY+EV+HQup2GLZ6s
rH8TwNLpCnebZu3S6ugk072CDjCs7S1QiVLTesE12UtgU+TJtwtT4v4X4UTiSnBiWycdMADK9zt6
mPWgm1IB63+L1rd3PxawQ7rW48kAAutBL2jP9pjoGmLvxrKgxhiFcJeAn6UMUIPx7ZwWVSnxEECO
fiQeYJpJyf4iSAq6GH53gXkQIVn1WhHJhpWKPZ3ng6JaNOtZO8z9FFLsHdj/lsjJ+Ww1Lm4A/c0a
toztDOP2FvE2R5dYJSvIIy6hS12SqUZiqzMoG75pfEB4ZQtVO13QMCUM1WMN89j4Z5OMh18bhC9f
25IXk/qaw1PCNyrW2utMuRdHGo/qodBoB9rU8wsiWJ2Q85ntdjx5hVHM5KYuxs+GyBM7CZ/SKjDD
R7qf0+kW34+ftrUVQfFRK2gt1MBHI1J0CZWO7H4lVIncp7M2iufImXd+s+BCx8rrm0/ZNW25u0oj
3cVQGJKIupoItzhKl85Z2RQg4U1JzftgusCqs9vCB4MC2Cs88uGfdJY06A98dzjkM9O7ThGl/K1f
bDLy/z0/Ixs/ionGypfBT6U105lxDqjZ2qv0BYZw1/nyZFJrDIuybhZBlhqkKknaIPxvfuPyfkBe
oquEvYLJrVZ0JMUoS0LUryq940YPdYK1h0BMc08LL13O1W/hvfSVJhfLJcGDHTlsN412aRc9ig1X
IJz3FJ+jfRD+EVAfXVietCOBTrSUMOr5Ae3JWFkifPR6GoxiHysmiJvR0GA2XP2nqd8r5VuKKQFS
ExmtJCT6ycitDCkzroTuqK4L4kWeou/9Wl7sRXCnwjchWs7IItwE2xH6tYm+bl0ybsvzweOZkT3X
cKrP6uyhvkmMrzGv8q3Dc8f7Kr+JEKBs8+nqxnwEs8BwGlKKEwZzLEhKFRBqK4YXuhNEb6isOgVo
dHMUiZJlKQW7xP+GqUOrmehtPwk/Vk3FaNn+G/swGZF6d046euhtQ271rdrQf+1v0wsr2t/WeMgM
AwH4FxW4HdjCGzQZ6r1V3OvWq3l+ZQ7c9fxzHVm6U1JU5CcbWkUNZMZcUu17N5/mw2ie9fh2TjRe
zxZGPmNy+gczqPslJ4ROUqmG08rbjKoigHJcLYcRyd1bgDyFPS4d6JAZj7sPbnYhyjgW0Nwyl4cY
Ma1U6oxIPmhr/y+ullgWlpZ9nDbyokzWwdCjAS0InIrtVgoSbtUqz1ihbhRchbjIBDsizTW9Imi6
BsNk/h5yreriWecfzimTM5D3z/KXXieA885HIIjl8f8W19nSAlmpAaUt6PFHjOObPHchWCCsQsDi
4Z7FEmm3liXA3kKHAUD1dGaoSgVKUelVAByKI/KZwi8i0Yb9c1t//XKatoX7/gIFqwl4GFxl405S
Q71bpcff2XR/OHVJJMABvS66Jwg/HfcP5Tf93FdEXQjLmS4wtBJP+c9V41XBkxM+mJvSErSRjdWI
47+aFp+ErBbFMMV1pLhHdZnz2ap3sMqRyz1eA89png694o7THoVodrz+lBN91ud6raMltlEAPLNX
DwdpABZSfLy68bfp7kCA8Ji8eRdeXjPzG/C2k0GrRX3B/3sIFTe0T7GV1/tH88dP4sa618fpLrUS
mcgJso+QGiGYcwEG28aSOlN4RgAfdsd4EGsB3hfTyCZEUpnGk2PtnjT5k+uF9B/tuOnf8tXNDEar
pKdxcw0hta/yjDjWNP4NSMkGvU7hPgKzxVew2xcAe8Izk2PS0Uj91uJa/mwhLDyThaJ1zbRcKl89
+Pcgp8GfLF8iCGhjC0SxorqgQx8yySbJOjetJacq4F6cfKQZVHhUGoTJuvzMdYo+6uqBY/JyG0Yz
Rwbx7pndu6n4jOCeY3NPaWLISPxd/3jW10HMGet30FEiFIeOzOPm4FhL4o/XLwGr4LsEfGo48aU4
IrhMN1V44TMbBmPccyhNGJzz9XaCRLoS4unkJXAheAyLAV/PNRVbTBjRiXwbFn9feRX+yqHVP9EK
CUgMIoTS8g4KrWaSqhIEWjINstiGzsyl45a5cXo33KN+gE1HWUiaFfOaFY2kO39PUYbAbapEQEff
uyw7LMvSd/I+CuksCGDWyV3hujImpoFZPx9aCdP63Cv4XLnhUaXDeeHFF4dX2caemfvi3Ah5I+B+
P93l9tGah1akeY6dlQMlo7h9/F1c1A4KruuyJOnXlLAS4zAUoPGwSUVUOfaLyZ2ng01HvcyMmSx2
REYKAqt/PeDymlo1x5I2C6W4OtHtWdWRWWI240i0lIrpPgJjOa0pCmyiFLD9WHH/9TsPFdZN6T86
wK1Hlh/EjwMDFaiiNa/0cJTby7A6Mq3anOGnqbJY6cXe03mz1r8VZtkHWzi8PbZFM/0ZTOBgoDfi
v4RQniH+vMLt40Oq+KNRcEhPtmFoaENzUpkpqKMR+Ul3f8p2tH1ziQ9PZSUpa9IqI6TMUjDIPbVj
x3HRvl4l0TsjkH1JqgVckjt2AtQmnpB6jpkJL0FXKwiVSgB2xbMuXQNySSKFVh6q6CdKRUwwyEwj
NS7Mw3435Yk37Ks/4+kwUdDMSOME3CkFBWoRRHwSB6jfcWzCiRPMarH5HaqClmGGwtl2CWNZ3quA
fEuqdV3pyVreMtqtic9XPf0Z33mXHkE9LU7l2p9Sq9Pb6CiOBzJlJNvAdZyq8ANEUO1UdbTSzh32
mk6gO/9kSSkkBtGtyxdpKk/HHnaTC6JZIEtnVuCd+cc3PdBq6ivYZqqYtqgl2SQIUF4HYSBxPYE5
VUB6lTeYC4JP80nCLzIavimHV/XklaEdoM4NJV3gkchLYQYNfhZSfHqIxxtWaIlndmQEPmJZUKLn
nKGuLTmUliEH+RT6Vc9Z/0dft0MHUSHwQVljXIH2PZ0TMTll5xoFOGjEIhuel2lecRWhgWsEFkj+
O8lr5jXwYOuE+fuxvhB+ZcyN0ORK9hX9ODwwb9ZDu2JT/gar7Xx5YBDuV20BFD0Rvh5g3UGiJ+FL
rx08QjwGb+PItJegrAQew+ymgrYNU0jCK+JXHAaxWZ3iK2jAmED56Ukh0ujd7C839ZHwTDkxpD7h
wgRrXHnWazgWEtd6IwOlSGiNeWgfIfcsF9tRzFrz9stzcDOR+PAza0I6lcOxngqDN/2AxjcBoHB2
+V1QC+ghuziEBZKtUQxGCa1kCO1DOCpmGWEUwlmWbcena4sKiAWVUlT97lG8gbpXb5cVq161FK+5
fIudZQU9XLqA0wfmWwoXS5y/C8zVOBV0BruiL3C1DZMcP4AmrhtJ1dBtL7fGdbRE37Wd1AAzaxxJ
7AlqPwGYVqem4sXRoiNP+v7q7tMqKwNdhg8TNckQmJDhtwNDMFxy/PBAYqeaGXqJQDsbRgrT49C1
C0qebkIo440TZoBlvgrxVimfVI51sc6EMaYh1VFZqjA8JuPSDydQed391IqTuV+6da9cCLgjGGqy
1bW6sD5gv0B1zHMPoKUu8/sJQRe+92FlnzKt3IZFm6jZ8kKcCyiiW1SBEgXJOpdrP74mWSdG3j26
cXk7VANysiPb3xBi31HMPSy7oDqkj/WecdKSBWgA8I8BnrjHinmPSPGF6wh5L8/1B2BQcFJmInVL
BCVQAU/hsba6qIKmu+XqE5K5xDyYzQ42EsYPh8f9WS+SfxANUIAAyoZaKDeQbsCNYUsk9DuSULQ4
G6uMsMmpzlRjpsIKMXcNJndnO0pH84/grfLYM/3Dq9Tt+0zQHQtE3WesQx2/56YAYOBM6qWLRw2F
hsXJDX3XfN1WpTeW/lFpQLDC472Uop8M0CroEomdDvNWD1FzEmkgSuhzf65UuVmMsvJNzsjT/JDN
zpXWzxyaDibal+OfHyXY7ExLb0TKRT2dZaYz6aq2NCW5zCqlCFIxrnWIMK4rvs1BJhETjoBc81AX
VwmlVD8e33zZIClDmjyIqQ4bYKBL+dRNpQp3A76bV/Vz7uANT94+UY7AVqSQkXLIqVoNb9dyGXrt
Gk7rFepZL03s8mK2fsijj++RAkP69+ck5mY9eHPaRGYcBfqhoU2vFskfzoQW5MgUuGYrrD0H20lX
DnS63j3hI01PQcS1QdIPc9f/GJtwG0W8ZJcZ31T/mDRbKTnWDaKMbSLXXkjaUq3Vx+O3EJbVc6f/
iCnITM/bbE6szY2CIs7avlLF9RGVZQ3LzKcfnMlINi2uQ03OEybUZSmHrIdIRZUNdglX0koFpYUW
7d0G1DYUPfy2hvNYG/JjNA+711vp3QKya5yE/vFuwxh1QhQWhHWiATc9GaYqMZ2Tn6RATArkO6j1
fo3OP6My9SjJ1Ci9sUcEWW+h5yErR9uwMHww7XxL6Fpx9LI94XwhFFv9SkGDQ4ffgmAyrnjqk0om
MiZGO8YppKKrozQVJQ/hgeyQhxR32ekxqOMaTovg9aYlqMp6VGUvxJPxmfjBLFqvD9wO2XIh+bcU
ZjX0PBOa2pPckPd7eMYJM3gc5yZytk6x23deF55C8q7GL45TESH5uAd5rpnWJ47W5rquB9vlpmMU
CcHMqSeqqqzFubJnzjlAnxbJbXbSFF3XhwB1+esLmbn5OXnxOHINuRtVx7ETWImoEUt24Hjkl9xl
tIc+rZBIq1+S7Q5Uz76WzjpFdTnM00dtpVP65ZcQnS+D2on4DIANs4syUuIcQBXbE2EwFAEPCUSw
uQrPdWCcKndHOf3IW8WtzZOyxGnlVmJ0ENu+J+h0IPwRtejI3RQICHmXlHh9qXJHm53cIbcqj+Pb
hZx+gLu7J1SvI0tSHup1XvRi3DK7gBC7K7fNnQQ9dlP24P1GQX9ioAKUBQNKB6+hbkjy5AIqBI4C
L4Tqe4nXFcx0EYxW3RmwXeI8NJAFrR2Cu2q1jIkKPKi5ZtZokkWDcitUaYyMLqasaWjNR5Bn3ZYV
1GHSMx/Y5+amcG/itLawNoy0A/FQ2RMlD6MG32nKXUqSS51Ygh16vRTaB5O/5DLRqqJr+4rHdnNl
RGsj6ncsS1km0tXscyUGvWy/D8NgXAoQ+eUl/IPFoAV9JUNSymwGpwH2KkkrbGRyt0Q13HYPv5dp
NCLeiAKoK1Gf4BXWqsJkU1jxeTg4dHbo8vWiLzXOPhqcDOeR3Yj9Qvjs794t9rwJnzWgHAaAUNMz
HEp5Fmtf7iAHb22TMjmFBjYWKvA6DUIdlJkPOQNOtqc4tlKphPSc0sar3h6AqSsvs6ArSuuj+L/p
c5lrS1MeaUWzSslnSzRU+dJcEaB3yl5zZLM/j9aVzmXGKDxlqfFHUj0K4sFxEUWHO5yWZVRh5B4/
7bHfuF70Lu5MJqkb0D+PLZ6P8rFed2gZU2Me+aVpZ5wcrLM6diqSatGuE0ul03Bfn68H64z7yD70
tX0JVki7g/TpzpLhFXHKlXX0a46eXUpothrF+AZDinChX7q0iYPzupwhLl1uo5+9RjbpCh8zdCSb
rXnklFzEvoHd2kLSRXyF73nyokKqNoFj8+WjAj8Ibv8PLSrql6sP+oNoZ3T4VWcoe116Tiab7Px3
BfNn2QurTwgS6wIyHCqf11bMdHKqisQHdZB9QdBAj0XeLdp5DrjB7sNx/lfeduyOIyenA2Rer8vW
hAhB75vgo0EffP2Lh8ItxlZ+ccVqK9AWH9nF/aw2bqekszigjlCu41F6inBPLI8IqLu4oVrzcNTQ
1lIT0betO2tg4rjW19Q7FjYzc+goZAm+bkge3/M96gXVIK1CGEgPgASL6DXN5bnxEtgjfqlmcww9
o+pgZeyZlR8SwojGNSWSJoceANcDbsD5MqmABSs7b4uj1OK0QzT+c2JT6lwTJne5S1CrEl3O8CyT
5HYNr7XuMuS5Y7V4hjt+IJj21zwAZhWy8TZk2bXBtu04gE7RXEHnT7paLWaIo0+uAB4gH82gtWyz
5EvdUcUkBsFQEzGlduNzHb7owcDL0hnXaeJOl/xlrHzz6q+uCBZXdwBxykKmgcOGxT2CJwOEuR5P
jEkTqV9Z7u5RX8vklAYNtSCjPpOzKne1Poy0muP0vpltReqHPfVmSl8SYtzVqoSbx6J+Z8QZAoYP
DUerUxN6io+Y7yepGguvRrly7LQit6JnFF4Fn2Q6Ssko7g4bHvTSRc+CiRkNvj1+fPdx9GI5Z0Wz
XXonck6HCcMfckBVslEDBy/BIvBI8m4iA27QP5wjG60yjYjDM6vCj5fviPvBtGG3rdttfO+e8/zg
4vAQBrxBpz4oOxkOUuE51hGhIDGDQQkU88P+f1isO5SCwgfG+tGH6rfNXYpbuET01VqMyui6b1KC
IYnGuxlKkIDbHH7eIaE9GvFB1elt4sYp5YStiaJcMjEpD2A2vY4njTQH2PHgHjwO/MN/KzfOZcKW
g5bTcApr05nDBUkIJucfVxTtRSJVyFi3XnBmoFUpFIHWG4lozDDB2lc6F3PDVatMzejS/25OcUEO
GZp+cY9uoKcCuUVw4nQwpAkZaaMeGgh7NC9AgZOCqNPyoOT5/onSZWP3YFwoYkxJ4J+5BBSkFnh6
WOBx3TWZvmVEYgfFWXj2+JEh0vCMiqr/8dlwf6vVLIkZVTxIiyqGacKkIfYop1mm2DkgdXrNxCnS
jhbCu+B7BbMTRm/33FqmAwSLiiOvRuzi9dtDTfq3z0DHHRNO7bGrbX44DHw9vuFooprZXgOAwacQ
cE5klpfrm3wjSrBBIWbFwnV7UKEp120yelmueQ2G45Y+fNk8zT5epEPQf+Fp7TduZgySZAPC3FMO
/MENNFq7aJmBO4i2WLt5sWgia5bW5TGbCCJK4iCoFfVc4IyRBwRegjQpxtYk9W/+7WWH3O1FX7u+
vUi+s1IAWMAwdj3IxDaAta87nHlMjfhwixs/j1AnVsHQIIoyLIQVSznnMcbKEsBeyUk3mR0yv+R2
7ngAc3FT3y98yXV/aMZLrJ/TKvAATXLPGe+6pjd0OJDYClyznJCGDcgR7/E4f+D8QSNAV1Pc2eNZ
qDcQJMlJkcDqB5UO1dCmOV6KdGLJoqpiUpIyzVb5Kf9lU2J0zYm0iWWkC83TA65MRTKCxcshiZo+
C5O90mjpyEG5p5e44dSWSOrCPy7jBkXH2SXbf1OwmV2AFtQKWHY8i+sXHlItPgTiJR+RJtiIemTk
spOjYFXQG5pVdOc477Dvu2IDyIhJWkugtZs701l6gfNWAH3Hrf3nQ1j5dkJfXIDe1Vu4opdUbAiP
Ocq6n92Py944jLA1cO44V4ayjN3ochLFMOB3KmYNWiiRMqJVzXl/ZTnRBNpJSdj6yBXvnQJtBKR1
zqV+v6tM+soDkPCSFrkCMu274SBT+T/lc/3Oa5DoVTn/tGTpe9AjIcAREVXJdY9G4jIptcMLzpG3
qVpSqQIps4XRrKse/mOeKj5tTo1lnEt4kwPcdfuwdP0XoqbZzRmvjRkPzZg9k8fVwbX9vBe7J72u
djpEttkIa3p4eenIiAx/EW4KH2g2ceUSULNIN88hqHPFkhTPO1gWj9Pj8hqvu5B+Ympc/yYMMT0h
aXRmd15FUqNOFEuF5qyqnfUK6r/4+LD/BXJiBnWaFZFqdPU5VIrBLl7RvZTs8XZNkMSEABS28nzj
7/0qAD5YW6fYaosTtJIti8LvIZtbHaPUvIG6g0uLjaYqsJyZEV5CX88BIMzJbydm0t16+5+I2Sot
Ikav122Z2m5KhMUEeicF9rqTFhsCSDKWc46xnhaZyAjxW0XB6eVRPA+SX+tNF4ftsTq8xen1Pbwk
X0WE6/z2Y1seBghUL+4S7vnAFWnAvu/IqaVOHkyOdgO/EAT16S1Pv5ZBIs2FqW5NcccKxI/UfHym
M0Ult2fZNNsNNSqxjiHWGxyKCjXLK1nC4DJNxZhWvk/WsB+VXNLl50xcIPEFNtHNI3z1ZFWtNccO
nhF2rLSkfWCzdJn5ngMuMbpyK9qL+sRJqPixlU67V14EZtwt+3Bag+1wIjrL0QRUb1eDDrmAABW2
yuFxnXWJufE9fySJ2lPKp3A8KQngUN5azy+S84zV1IJ43vX4uScDPr50TeQFeUJCDblSmmH53f1b
egsxNTSnSXCyL5hiP9RLYUkD+Doar8W6xG4KnrCggrn4c4GFrXDLfkjapnOaYvL04usZK1OhawUd
VZiZ6m+IiNm0QrltlCP2VOuF1ByWq15P2pQA5/fXDkt7dXR3rQeLPWRuTwv3dlQTx2HNQw/bPCHo
gOXM256n9dbEcrALc3+CWdCH8HFMXU/p7mO3gprrIBxdB+FNVG7P5LuH/pHscXsCF37aNX+8dstK
QDV1w5qJtw90YO5p8Ohtpwhqgb583S7QE++oWbgweFYTod5FoOqQujgip1sOGjNY4t8p976u8ouS
8tlXDrmvgOT/wXgDBd08BDMol+/MMxqgY+TmjLCaByWuuXTyp8G42wS+nn9U5/Utgf7zuJdPRsHc
+++nFVRb/tWt4s0fcKfrpl5bAz9W9TpuiWqselqXBp7SAIckRU4P0hWw5IptzJyjyhNl7/D2uFQU
9CbDM9nAwtxKGw6+Km638sCNO8ontTQD6gFflofY4Ww6xL6NUo2JsldD1F2xb5dFiKyyL+LgrFgF
eqW2IeYuSEH01Lwy1xrH7f+A5hFx16jjt5EP+rkA/2uX1/YtIBceUHjsXmdSS+OK5JUfmmG3N9ho
C10S3vi6pUXHGlj1nBbwM6Wh1mKdafi9MvbhjmfisTZkhQseCo7ULKk6/pBSuCLZBrsVKoF4R/wv
/Xc4PK5LCDarq2NbBNmN62WBGkGDBishkGt8q9+iTy6KUoeLbXFYkV6Gw4ewCTEZFVF2dSbOjJky
GtyKfLuv/q1nARv1vEaeAfqwV9dfArawbYDdvrP5baE1V3hk9sVdlmJ4mt7+JMrjTyoL384VWoJP
Jm/R5IoUF81boTWikBQ71YalekNadBpJNXYv6LtAo0eSrT5f5lIGgNdBCIpCi7dUYERMuYRn5WGU
YFhubv7h+112SQkRbK20Jn00iH+8GYmHK2QFiH9yJGC6DEOunKjlq/r+FnCRFI8VPOAkSU1PKf7x
TWj3kl0h5KJjkClDcWYjaAj5HgUYtoLtgyUiXFw3VV304346BUGcJymdIfukvQyqH6Lomwhjqbs6
gn0KtAVUKnEH5FawClrYsNHGDm5dE1YKA16/MT8s6QaXXgM6NF0Redejd3duwbjSonJUxRG4DmeA
N/XFINVS7yGe8YymaagmCVQH/sZD28u8BSr2PerH7oiseBPbV0veNq3jqGDgYkuwLzvt1xGuwOYV
4B/E+DrHcMP5HD50dgCt/gxWJmXp4TbXPX1j+VwNRcZyDDMjJH8aKWn3/7vwV3gm3spfOA9wGr6A
M1MHXY9GXbkrG3wu0Su7KsqnGBQ1ioW4BZEyM2gvOPH9HfqqfXAMAt8DUqVOCdwTobuBPzuVcKnJ
8Ldb/YhHFx84clBgwyJhlcnj1kDlk+5udT+tAlGKISRvC0CQWshWr1EV8vdZozuQFsrguK6/UjXO
r9AOHCIOeE62FFVWEE4iLPj6dMrAH4hMYV98KDlHQx4XiDGii98vcOR9gtmixrAgR7WyuI0sLcFb
Tb7jx6zHYleGIiVTTNsQl8oLFypqYIv2lxSt7dLFsXxO9wIDOMg6/UAdUvevVM2mX4UU4/B1rZ6h
VUFdn5F6N9EziwAioTi9CWL6RsZboKIeTsyg8zzayFjoeU9fEpvbtRNaa54eQY7bKYxOBnMrijFN
MpKmLDZNITxn0MwChoJ6+h1NNNl+NeGNlkRUDalQW2p4mtSeunGkIUc2UWybhWGB7/NWU4pHVLA4
McVdatWaw2GOUuFji4u27sfmf/OtGlZF9ZGh0XslwSdS4sYwcujAkeGnshWwY8hHcxh+rdSo/VQD
4ILdpeEGLZAQFerJuyVBM37MLn8Hf/wJcJpfFnFAzq83RlpRLRhJRBff6aOqizY4EQXBTl2v1KkQ
1rUJKedW4xmK+6snGH8/9M0bzGRjt0yyLrsFcDxxHwHT7xeDyW2/4TS4XRlWpq/pgxxiYogNDcUs
lFBnuJV0hdjSusLB5yIcdXAfkvsvcIaTEEZRo0aJux02jz8IQi3dnKHe716hooNv++yE/pBJeW2L
hnC4HsPRHmBhylaIWmB5bP2vdmQa3jBMhTfqRHxbpWnK+P+H2inUU9ZmlgCwtFUSYOWMO5ED968Y
X8PAJ0AW6ZdUxN6GkAKFvnKV4hWNJgFtWT6wPR/7bpZq1lxAQjuSCulWZ3PIZO6q2q8hXEMrA1cN
OOTM//nLT02ajRP3mKqFWkQ0gS+X+oKfA5qVGorBMT5WF+hItjXjRSjoat5OGPvxbkdm8E/e71rX
rM4sjRuTA3f6JgOdIZZAaR/UAn74BmtQ77l3qUNKBU3a5ZQqtw6kXlN96HIOUf3iDsuPTZ4QLgaJ
X6ITvi+VctA3bde5Qh9reoo1ThvF4faS2HOg4o55TuXORsMqpU3dRfvVTIyIdVGWfmuKVq4OIqPD
XCk6+du2b/SwA5VH9F0b2qJfaDCTL1sbL5cvnsLFw89scmGt2WEO3M4UQVtDwIO5Egob4EA50T4B
hc0i3gWlgplDB0sf8vt3MyI443D4fmUmOQfK8cs12zCxejnilRAye8Es9tRzyB/JSJER75uVWsp5
anotU6MjWXwj4/75t1PNmFAZ0DN9Th6prRIgDBUdGBmAQGq66O/C1cLY31bFQX4F+AFM8ZLw/QQ/
StPnd8ecJGTHPUf2LBJsAbbJnVc+X4tiUh/31F1IbwZi+bxdoZGCdkdjNo95MDLG2oHxG2wbBDLr
rO05Sdp/eM7p7+0l7jmMN/kbiS/5RcnGyHqGWXZXW8eg3kQuggLa8xOUm0uaVw6oDHwreaSmtWFs
ZhfxWfBI2r5pczzs54FxNxfFz2d+SDGH8obaeoaZ05kD/batKTx1Q87GxFytce2HpB/6O7M1m9oP
4whYtQhRDOlCjFCzcPngqeP5HO8pyjei10qBKLfEm2CAUHXTOAi9kYwG/iQjGnetPGKrwWyU+/K9
FUIRf3XfHl0YpLUbTZrOKfBAF8AlzRHdLk+uHFaglZe4FEVVoBb5ARjq6Qb/zT6kYQF3mg5D2RzT
XioaWxOidxHpj0u0X5INsEzjq6QRPPQ+8MbPjqgaOAJcLDYRNbpgqLATyAvkUmvNZXQ4JqEJdr1s
SdTj9iApYFDqo7+pmAuEPLYPR5l6i49H81LdRdLwMk7U2YbPrA8tL/VJul9Wv5cZvfqRLZbWi2aW
syMEq5hzO8RdpH8lrQcG5u7F9INl20L1Aup548jcHS6PG/k5yE0AR4JNFgcGsEWbw9WrH7cnapV3
J66GMUVP18wnwk9hIsWLMMYNPNxZKd0kqUA+Lf0nKl0ZIVsheTsmMLYM/uavwk9mpF2ZrJ6kc7ZB
SmEvmCoOhpVHCHlgclyrv6aImVwuvti1INndlj0RKS0RT/rTC3P00BW3j5IZKXJ+MSU/Wts4mafn
1dsdmwLq4pP95xVmFRTB4lPrL+75NkaH0YlwQx93KUgDfvGg65Ac7j+uG3Cv6vTa//Zll+nshvLq
LS6qemuj3zLZWs5nIRLvJx/EKpBQawsCmwPbKi+bzVcR3hoQh74cAXGnvheC58qRcTw8A+wgv6DH
6UFiu9FP+jsXkBiCDo1p3iZnNP3YRiXxnpa97HhUBNGpeyMWPuAMe2OOQGup6ta0/bwA0A5fDtsA
JbmgJjDb+gf3J+9rtI0QF1w15ET9hIza/ueJ2PAGimFJ78RUcqjD4ZqaPDTMxmX+aNgZ9KYs5a+V
DF3JHgK261FrA+rk9V04NwotQpGK/ecweqf3eEHOcPsjP/p3MltCCzmxEmCLCx/JDfykPoVBZHnl
WVjPoQVXbqHi8ul/pZdyrEKgMKhR6cC0J796LXIbBhZWbDUxp4tNDWqw39+CeIaC2nVNwt3kjZnc
WzuJsKLfMgVkiDAalLVpOm4Yes9uRcNs+/gIYMWT+gPF0F7HyIYQF4Cs+pD9OI5vonrAkqaAoQho
MM9+q9voBF1kPjIHMluU/SiLQ1dQxxKbVHYlaiz14iOdBGmBnHT/2Cvj4a7viGjCUVln/fQ7JNxh
AWViBqFkXVsxiGUpoauVU7nKOZ2J5CRNkAeGcYeiWCzNufuP+YMmTIbBcWQeJ14fuPWBRnOhzPTQ
XH8wDN9v3nB5mrDKyZ5u0VX3pQ+J5xUschruFCDVoQdNWYfuV+ENjiyajGstfrSPb3W3w4qBg34S
6SW9o1fc2G1/Cwr1VVHGrG6OA9I9ngCbqKukMXhJ9msK3J7ZZlhYS5zrdWfBWZpp2mrQAWL5848w
G55hKujxTljZMPYgrS91B6pOVXfOHxO3lADhNFK4xGpOOjDYiHyNCguFmLE8L/KfuPeWi21C82+q
qi4z+3hCREXkYha1eOSu4gIJb2saqqmICgeKHhad+J5Vp3hKhcSO1sB3MGynPnRtEqRYY5Aw9jKM
MtRIvm+zngEhIsTfram4RL5WyPK3QH9Ydd/XzP9iURqXU8ImMeHZJF+V2bht1FPKg1Ugkl2wq7D5
g4KC/o5gbeDg+z9bhxi+5jZlcqbf+Botf0N44wEBUB/pY+LXXqT2q4BWxnDAkuXJQ7P6XmvAvXhm
H8H0Hea1rzYBW1wjOOR/mWJYP3DcmVOFCk/LXZfsDxm19hk58qvCP90PdhsECiZPPqqptJ/G1KiI
PtWgEgEcvQrm5Z2FnZviMxZQCrZnIe8k4w7VGoCgqCOGJpyGjWWiVpHbB/p1KyKQ7zNLaIaGV3lL
2djh6BUe99OMkTO01fd6qfggpdEiGoQnFX82CxkYtcUh6sr0SeE03dFcdQWJIezzSixjZXzq5HKx
CW8Ru7OPUJmza7cm+4fsgGa7vUJDLQyGWDVw82BUf1/snOSVGAkxZS5lDNCgVugcoXy+SbDJXXEf
PTjUL0yvxL5oHOSCWzvoT5I2ReyfAYJyUKybWUbkAj96AnKAjZodPnFdzzcn5lB/MA0NOUx4QVx6
EVqYY6qnmI8Q2TmLP9aXkElZBc0u5kRRqN8CD5fHBT5N4Z6rJLjEDP7qUr3LyuYmOMyaTeV2r4YQ
z2g4zvLycVW9669w1O3WXkgNST/42xPEmcDFAgXMm5ZBF7tl6MelG6gYGa510BPJHb5xupiWLnsU
b2mVU2aPml8KHK51MItJ459L19OpEga6v5TpznD6irBDYu0RPiRyDWtH/9VU1QB5UBoD9dd1P4Vs
TT6mVPGoxxRProS1dvRcc3Ier9QIEFMXmSC49Zz9Gp1RFqsVtdZea8TbO6VUu3uyXd1zbZ8DUMmg
mlmRO3Bl/asXYniI8euV6IxpGrpl7X9z+qKzssfdgLM1f3AMLTjmLh7nx2F0tvh3r9Uz2EYicE//
wx1oVOY1bW4LziPp7gkEoO/pEssLSC3WxefZsZSh+zjfhIBfIv2dk0fkFGvBPG2LshAiruZ4sFhI
pPwU3MQeZxz+eEfit7f1ALcpi2bo7A0UUT/lpYFbdD0TLrSIxJfpaXDG6MQj0miRRaRXkoA7PN8G
A2mOZyx4/4DRgN9ZfcytBxpJ8Ou4hKu27euhhtaf2la4xDtUdW5CLJncFnTESCJdlTiW0nO+cmyw
l4K1oNT4dPAsgvoDOW561MtqeH28hCLOLLg0FvGZKaCIFLkQ/wrJJUGaGur2UkwcB9j+vTiYPJtb
nPo+l8HTwIxr+jyWO3aRBubC7Jp3/GhuG/7+qfI3d9DkvWJxTGwv1PFUkwoVKcyIaXHUvOy9tH2r
cgJFbLZjLTHatuTVOFCTIrYTocVJVzu2PDYzxoiSRb2KT30gy1IwCHxN8Y1q/IsY8CY0DTaKXpU8
ph4Gz7pP81w8g8mmrUDz8sHCPg+6eF2ONTpLTbqtzMZ/8DSOyXbthq8vPI0r/o03+zLEDoTs3pGE
S8bvJCFP3V28O7eqS2IWcqNWc2jSAuuJgbtiLy+YXForWGqsbxG6FAsr9skQOz2bN4F2fmeN8U9x
bqM+GGUxEw9b9WTsxe1WBZqxy5xLHzF4zyPQZxlv7rozhjkJRWdZj7YGXT2V/WhdaO53Qpv/+yoI
zBUvHMygfVmZhXqD+l8a0OazgP/ZUbXhwkxgOx4ds5aOHamwR4il80F8cfBSSRFbghzlBk1oup7e
m4e0YxfRpw034PlAjktlnDA04u2p051FCq4FPmd1VcS9EK3IUG7p73Wjwe8KZZuwDXRxXBgjDzMw
mqIA3iEn4poKasCfk+xIkRPnlujkn+gTmLsFRt7vsZd5XtC1hUl5K+xAQRwbsJhK9Zw3vdZ1LmZR
ErCqgWGkGPN2BMGmDL0Z/PBIBiXaxh75ulADHWwV4VTdPiNSGJd/CrJjX1hT0Gq+XL1q1tO1rgSN
2RujLWOiTn63G3gYovILgKRbggEdKCVgbfmSb/tJZNmMZokvj8he8OvOJA5T1W5UeGb8F/PkijmW
bOOVYxOFNOJ9Ym872bCJ8uTYNvA0NVjnhEu47zGuOdbK0gLczaB3YgH2HsxS0yRZU4YVP+LCYHHd
NfSNvIhA5sRxHHPtmJqjrI90RXMgdGm22CJIPcXko/TyyH700sRzlnlsgk4Uz5apIbx35Y/oijjF
K4bMLrriTwerC31pUU8BFlAFzSE53jSVA80krXpoRvHc4GZs1/Li1qZ7hA4R9NFVXOCX1/Jmf/0Q
42Y687mWCNAKdjNUW7AjdSIfYl2bJdDV2mu7wPekFS/EgogXxXmMKvrHK4dfYvHRcIzwpI6zykus
ZMGdLRM2/51L3LFDI0PV7CFuYt3rRa3XW/qudD/DclnrslivIsO/UQV2QNO92+0wN7U+UzE1bIp5
MLgf+wTedJI+kQtrQa1JeLfHMDKvg1ZXq2s/cxmKJjPTrTn9C2khQ2S/7bt27VfWUVdHh6uXYoO9
3jw+7a4Dsn/AlH8MuiIVJ8PkuoO5Y+P1HqUm8/3ppICdHTuyVy5DWse4Kt37TnRrPhlP3xUFanlD
+ZAUhJx+0HsvBcGFyCCzzOr1bZ91q7MjSbXLUuFh8te2/zkw47+7YvNLJCThJUq0HgJAlg3AVOcW
GOrGb6UQ/hfqjkD/d1yQ99gzOg3/XV6DizeUNxkQ/sOWGqMuvcA5iiTPEhTZzDhQ5BCKCxtnh9Lu
mtJXSrrdon2DPEb3SQqARNa9KbxHGPun9qwmjeZZX6D2FlJ32+PfBrI+mJnsCKpLKivjX4ATz7wU
tagX2TEm7fNZHBNYpzihsbTL6ieeex54YMi47tJlNf6WIfVjmg4g9d4MYeOetr4iqGjaZzbmoZRE
Bnw7rsTAXMhC7mu5E/zA9yXW9t91wvD2qhDHKnTAMtWfimKKjLgIMUrXfkrCcYrkpOeK+uy+9y9p
bxY83g3FMugrQRO2f+W9cMuBPJYnYu/tL9A3RB1oGAcL0sVCZ4hlbv5gr0A52S1NEHOVRZH86MI/
XyEULQWCiJBNrhmd8yrRpA7vWOEe471/PCCuJ6o66kFSfbJwe3ToXCX5Md1hrGlYrygIQ1A8BSHk
KqKCPdj5qhO2XG3L89NjcXV9NtDc0354P52Z0x3L0R7SZ+KO8kG0bgC4ttA9At7OBhAAWEqsVc6D
7s/Kk1rnVSQABkoUndwH4h1aZ7OtPpr4acf00IpjKKb5YmmZAoO9dzRCLrMix2BUOCzh51yglhAR
ijjyEaLFot0T1/I3hfSUlvk0B+s3TsODh1rWoJ5ddYiFBG5HJTglaWyKcTHpF1hKnr2NabQKV4UB
XHW1O+Ttwb0Ao/xxO02JhQGA5qGLKB7mC/59FKxYQNI1HyY0R+oEAA8Ivhl3B8JUKNpd6IeTQGq4
++h8VNc8jW83Kzc7iv9eRB8IjjOAKe8XTSsBREQF2gmkkEqNv/hhCShlTUAQ94yXetKvusYU0uEf
9JC+AEGTdgxGUEKQfRibLq6NHRjIAr64n3ebPm0GhOBh3FTwG9JNxtXb+LQGCXQy2C2wSw1VDpMw
i9EnfLzvQiAUB/UfokWjRN8c3FibBwueih33kHjKyjNitWS84TbtlsiTg+cK0mI2Pff3bIAGogrL
KdnUQKGVE+umzj9nnx9ZnJeLZJzQWJzjPVq1Oz7CCO+SavDMyqk+tZt+xjgoakX6lUBDiYvTyqn8
/GqhnYaijrTOY2XoptBL/tMro/pVA2pYKlW/S1tm7gsHgnx4LRuMQQXsnxVOWEubuIJKSj1KhuaI
nusttQR3hP2mMNs0IEbS/X7FCxEr5Avi20Gk+K68YocbVR1DnXXef6i8IvAeVmAZJfbbJsdwTEiY
56cjguySXKhVtfYFagiZy5GKJuaEn+2XfUDo0EdES6IBQ0VGIXGrQvA88tROmsVMqFIaR50iJf1b
sb5uJO3E5AdXgUfG4mKQNVV8yGlETcfGRKmlrL5F76Us5Z1OrjFE8Z9sIh0kaV/p6QLD5Rjn6S/A
s+GoNLwmGVucXz7VUzpnUxf6p80XxC9aRp38g89RoItag9dCwB+749GZBD0Ju1qm1rIL9gt/xe7z
/rT61vBCoRCvoxq6sE8FLZcNyBrNpnHsQCZg9Gpbs/MZ/hCwWvnxTGHb5BRri1BtfLHXEdR4DTik
/twY5qTd9ZGM08Li+rjDTfxsLxTznS27SvQAilfFiCLd58CrVXJ3h8t2ODO+L46i+kSNDe4zp68C
hDsm46OcwGyafRhG5FNzJwYEcG2IhhN/DhY4pf5NcV5ITlPdbc0kB1F5LwL1dAQZorsGRWAbwKkS
EtJ61x2qgPEuiIoRNbIAZsbbvV3g5y8Lg4+3gsy8m/marYA2czJYf0ID2daYOrushwxY2fIuyeP5
3i/sFT3Uu2yRBGBblsv+eqI1Slb0Q2PRyfm7JazmLDEOlh1OHKiujGFOwjry4rZXUEDuqRLRewNS
H6Ng3Y3+5QgRM5a8fqcmbi6vO29z5MOm+F0e7dg62QBNwzNdRk0BNU8TbCZVtzaoGeRI3Ndv5upn
17h1/+xUMPZl/phdiHgk9phrhwA3uMYKWw5jm4E6SLtfaEGda1TJQn+ZYFics2SBOEHDw8LGkXdb
Npfknn9yCA1H73Bchl4XTwG6SJUsQ5TL11pf98MYpN+ksBFBoNKOCLNGIZxoQQzo5j9SRTwZZ5hg
vCIZBVypASjnpxu57mT8KJ8Wr/4N0NofkpQnd0CSgAc5ZlLJYldAkEotbrw/wTZcv9ncve2LaEwW
AusVHsFsSKVHwYfYaIMmgneTdlbb5lJK2RePc4y3bCds1/XCNd0VOuOZSp5I21ff2qyy3O2Ys+yZ
RfptTTmirsg1IF+eYnOX1N1KMw+q7K9qwKB7aMV9wnySfpRmN115L7A/nUc4cvXmRB42dfuhKpYF
LEKNSeoVBN1l00nZhvDVLdCtX7q1LzN9PHy8TN0ueba/rBkQPIHogLqtYTTVrZSCXm2uH0sXnhr5
2EY3SyVKRgv1sPJN3Gq5LihLZJAxDIqEtuzwx3sgHAqVtNuDkk2Le15IQ04+mFhiwsdRn84IiXJi
Jd1jMVsEXc837Myut5AQxgIOOlIHaTRbZOfp3adw60UjfgTx58hCmy5cVksHSbTRsK9jb1ITMTvW
spqzDq3IouugEpAsoRvg2matfnhyEi805oSJC+u0EKt84iGMalzLpOgjMH7Z9eGoD04Z3cDhXrgo
q5nvIWmuC9ebrrRAjAfLhA3dQTk7N7d+kFGB/tJe42onj8qk5dvwBaAhSoocXtRfh457/9iLmJWp
CuIlmy/fXu4xqrv/AmDoSWBB94Njh5dhZZBB8vARn2LWax/6m1C3Ubvg1V6zogcnGzSOtA6btF2M
NuP02hv6sECuIQ7DI7uCZNOWSNLedKENECRCR3LOr9utvO1ggUNhiE1a7ZG5i0PxEfAuMMco8BAo
QS2QvII2ni87RV6V8F5ktZdeQuGGR/WWBfxrfeYEAUeYRk5K57c1FWfHwKefLNvCUzdlNVew04a1
lkwjWOlsQSO/iWTOsTEQlxX4H6LxmGxuDtfLXWY44aQ4Xz91jfP6uUN4ZoAthTaQdW1Tho4HbYO4
RAS/QZ9siAuQnjfhnImYKGIm9eaygX4Cy7fW1WNUBKb85Ay0sG5iHzvOr6OSaBTwfOiVf5YEO4Jr
Y4XG9fjCpFmz1pFvOdnfryOQMSVBNWOrTzbH72V4oE2lG+3B6RuUE60LyOdN3y81jDQZng1ZOdxO
9QQu70FLVhFIFtpIrjS503+7VpVv0zoB01xeO6L1NQ+sqnA17mtjbqfk+wvsIUvxspwCiXb9HdX3
pySUIjsofkAuMELqMnUXQfZKl6JCSBK/sAwJiAJSKEHOjFsOVILIIYTxnMAcx1Vdb+GShz2+0NPM
1XqRJ+CZf/uicwmrH+ZKPc435+1vZjt44ekYwn6pU98QB2ITgsGSd0epsm8QR0uK9/xLpLvxIdJd
oB/gKJ+2IdQtYOVYr7WbaQuzxAOvNqHSGIcLqFh5K3U3gAgHFC4tyAtDeCFi1omG3MHfzvdvmvf3
HD692Cj6k+xw+o0Bhi/3pf8GdRPn/G5mwVL7/oQR0qDEerDT0smK7Pi3q/xU+//TVDiVkINMZsit
vQaVKGxptw5r7QRGrsVYdI8vdQKwzy55ieuOs1aV30ZOtNSrCAFAi2r9Xidide2t9desI6hYGhsD
ZB91ndNtmEz3o1hxV0DwawOTts7rfj/rORvWHtRSPYY1pcxpXhQXpUGDesMdBeP/wGICHbDkICNU
TVCdOFmXzBGXPsX1NWu5Fq/JiIUHqTFL1679y3CtWIS4okv3UwYbJzO1sKG/VNEiQiSK3JmrtvSm
dz4S5ua4KRJ2KONvfFDzB4DbLEFn89saETxrrRx0AqzVHGKMLHUojBNTs3RuW1/ngFuCGkstnkVd
I/SvKXjp3fnh0V6+BGcqLDFRQaFrLIOvQ0JCSy1PhV3OpLP0ok6QXeQsSiKPQCmL9GPd05OpjCKz
hDxBl/7j6sPHHUEnr6JCm18Qy0R7uJ1ZejdQZWA15tdZhRa2XKhufthSOEwQhpP/5jzrxK5hfiTj
k+ZWyhNbEFRcre9QmoMqNSmGq855Bv5sQCcfCbChi6rv5lTu4fNGZJMap91/my851V3tf2jIGnt3
OT3vtcKeisXvjsRHOIdGS0wYT3po3lH4rG17bFDyPbKSBUrUSxrzh1j4NXdhA8AI/a22ceOfHwzN
DJTNm40jDzu7qtNaFC0J70kHneT6B5DnzaqAduH6t05ATDa7oEb9yKAg+U+VixLE4wMACpwKvVXU
ZAEpyM4ll1St0urAD/Y5rBCKSXtJSHTsqWJD1sqQ/nRtArkxWa/tahtQRQfrJl991tJT49NHaWlf
kFSxhaMqKDtsMMKtHmQf4u0tKOYi8z7UdC3ggOKrdSeG0LTjc+eF30m2YYdxtproM7nZ0ikJ+O/q
1LAMg1tL3Ka8FSZ7jrRCG4TX15huZC7HwjMPDMFDL2O+mXDlyqJGPxffUmKh12Eu/tcw4OSl2TIw
//FDTnW71891/5uXpHpDqwzD8lsvdhYLhNQ8fRXBJwQhTF7a90If3BQ0Bx079FfKxbtRhUGTUDVp
QvMs8eS6Bhi82QayYsz8NXZ1kAhY9Nxr/2RoyWEAdUqSnBFMPi3wZD4yQ/FaEIQoSY4RTPMP/X+x
hRYVwxvYsJ36Tsrh7EqP1IQkonoSHucf/194GMSFS7TxpHKRFv8+aLr4pUfmOafvyBYwKvWgmr4+
+9fcnVMqVbg1gU5UBCwBV52AbCtrNSRWlJjt9IVdqHknalTp/RptJKSEMb4rPcZulE/WgwKbEAYE
8Wi/Bei1FRxnJAY9g7YBJ76wJXmMYFnw1Yapy5S2jlP1Vfvc5YZV4QKD3o8zEpGTJbIQC16v6DEm
jPC1UgDAzIL8FlygEf8eIsTFnpBm13xsSFr7xWALbmswK8X+9c0YhSNtciZpEseohnEzUO5mMfog
GgDLIp/xrAbTrd2Hy++i3PT9FVJ0m1MmbsBtArwOLURFB+RpyqeYHlR+JZC3JQzz1V8/22oRDNij
lAvm9TEF4YP9QO7q+Xs8/EaM3OOoC5/Yvsg0p0gohUijrM/yzPsJB3KUVBvmCYNl4+5qvdacIgop
t5fOSUDJvIh+UPa+E2e1NAbhc7N039bmL++kU9Qrv5PzjeCeEnq6Z1bIFKH3w6M8JcBPla8XLGiH
fl5sOK6XyEVzRa0tySSYCUZ7TQlAHFRWPtjydEszidXYStewY1/InJekj8Bw2OxVsqC8p14ikQyP
i4ZovXzKhxaK4xMvwc3+LyLkO+qut/doHjaYGTqDuJQ0lQN6STsISF1DErrYb62yEWsfZnAbg+eN
oqKOIy3Mc+6z//KE2uJf/hOZXOw8uZvdJAfRraeSGiqddXIrspLsiF3Bx3oY1OelDOEw3Zhc5NgW
Wi/I2m3wEKePvLi/5OOcz3kEaknZQfWPCgsTOEGIVWHlyHtoeaUP75X/8l454pS/jDfuqeTvupDA
Rb4mS6X0M6YGNlYVsvT5i2NHWesYAbqOsMpbZr8NfstS677xmbnA9B1FrdzzWw66brH/p4jsKsLZ
hW05G2LqeXT9Bocfvaza/Sq+WFvyX0eHTg5A4uYF+a/XVIkybxLT0muEJKUM7RKDzCRn+SdYqLAW
QiIiyrqYe1W3LEE+T4+pkVIZQrJFXWpHhsAbokjmFZVmlZikcU4q+RA+P9JvLT/8JgcehM8Y1fMw
o/3lHRvALDkuQcF2HCEtuQITWaJJLPAz7H6x0Iwa0Gx8lHhle+kSgLelCF4t9W0tDqsEYeMhe0UD
va40I/hhUhwe8xlB644SGDWGJ4OSeHs8unSqFD05PTJvPprdl9g++GnYbDeWgR/35MxwHHPs/E7k
fi04TCWZS4DgVwfQwFsV52xfDcXAEJXroGlmJCAYdfeH+LwVQkd76+rCzP6sdqqc/emFtP+7ldmj
isAKFed7uWwqbBsSSAazsoJxHuN107XueB4S/wBrdixKqfP9J2C7jsJXLh/osLKFXJcBAbW0CkeM
e0JhMHdu8J5CSfDuMgLz+xvj0FH8YNZ7GhEy0sKisalh07ytH1rcV/gEzbI8KbY6fOHONc9OF7Lv
29k4owyjBt90+16AneRUIUqeAcC65x9W3FpdnNZ87ppzLLafcS0fDgSClCsRDNJvptwOeYeSn78F
4e6nj8kty9ZS3DvHb4RPJjRB6JrdtPVOpBU9jGXEHcC0REm813ucP3NKRd3YBXWpLTKqjw9trXZ+
lZR2YaCoAVKHjXuEgvQ2njGVfbeWzL/B2cfLKBO3nKjZrBUBXx7RmGQ50PAlvEjmB0HUPjqr83p+
oz+rtjjjbkvRbijobXqpTqdYNV/bQesPzHZuWD1BNxOS7uOprjlql4LKLyhnpMVzi4pBBpubivbh
9CcJ+zBQeBHBJ5o0oeG3XKeMtMDuqd+ef7Eika/vQVoIeK9y2Pv+w9YBvvYMcqtZyyhca7FlWlgq
PmV8GJwNIkH00g35b61t4tLJpsuy0UujcE45qrT//uOwI3OJ5LzxGIzf3zyMSAmTWpXqrvrSeZQI
ToaisgpROC/AoK7qixSXkeGWyIkxzioeDEoZWt3bQ9r9gZuuBueYeP6xELmjirtmyoYjvV/o5Pk0
xHO0OMfUsVmVvNlDMz66D1JFpygWLtXwYMBPMy7MYiiq+CqpeDIOMMggH4VZOtbP4W1jLteUyYoY
stPJOTOFPck/ZaZq81CibNtz5MxjK2siLbF9qI8h/c+J63Y3Ns+67FLhIxYgJOCa/Tlp+ZeKyS8Q
61LKUN7/ZV8xXoLiOuAcbwXwfRsE5238CbTMTCwN0+da61Wi9qXFWhgXfuvpVhyxKD3yWDPQySmx
VlBfnN9CYeFO9DD9bnDWJbDNb1PHuilyB/lZEFcFprSYh+JGyk7QDjxMbmseCg1NlkIdJPCFu24j
qa3n04YT/I+siJGDMHIZVORhaw8guHLksCHAZ6/g6ydel25BVeXpNL5fF3nL9BkImzuZ4ma/L0yq
j+u7LOEwW7ykDb6GuqTD+/MOwdB9EYER26M3F3JGaKkBMB0algvrx4azq7nJ9zEstDuAOS8oNCHg
qzxxD399XvXFWFLAwTZk0dgvA9xUDXgVHdRWy4KhUv2TSArERW0eivF3EJclzo88DVtjYPxsq++A
QgsvdDJV8/g6pcji3MRVMCM4+PfpQV7gNDKUsrcJs+4S92rl95zkGyNHGG978wuXowF2aRW6am0p
sl+Xwha/LnfdxusBp9EF1Sq9cFin3HxxDABVqdtAreKVgfCzXqda7t0EAhtsM/1/JlPPcR0piV38
pt5R2ELEa+W2+wfrKQ7PQ11juR5Xs7O3bsgs7UzHez7/mdBYXqiV9aqyMgLtiTA1xG6CA9Vt9wnI
z8CuewhYFhd7L56WHqFwmS1W4FC0VPiJkHFFj+E8RZYn2YjoDdwQi1jU3U04UiKLRxpffEyEyvvb
VsPVhZwkl08qHmUMXFfi/K6eS3Fypbtk8G3rkzad3Cm3tG9vDbo037nZJu3+ad4nis7g8mJR4fBe
u5MNTbYsVPhM9/aPDC+xgZlJXwTQw0MjTD2pnrMGS2fwTAUhd+qdr3nWZHzXw/1T38xFtUTlscJU
wbbRNS1OVTiHfkJMMfT0QMTPu31XXgJCkfL9ah2meLeDkZwMngVjosU/Syxl0OVWerfJUEhT2Ofi
YeGPPQVUfeTdOmlRGbmH6U3O9FmqH5yDbTBUqO2G3vj/zfsvvoPQRSChuhUzIj07OZjjPtW81vyC
QuLutYh8M8r4ASFXJ6ihkLGRbwE4IZpT05Sd6Uo5FULUWpqXqpLKQQO9T+XEca+BfjXJpLxUcQJP
3EPjEE+jUtuAZfdnz7/GeIlIt9rEbGRpn/YLDk0yVxm3dWft6NNZJaF18YW08GgkD/xYOZjhYJvH
cNsP9QJk9UUXk5FWp/IDMvlJnq/TNs+lTLR5C6lECITr6UEkElI8KNup78XCvzDEQibBmQxYJtQI
WCsZ6IbKMgrDEQOoGHuAOkQxkMBWPyBv/sAQMmtvkZhJ6wnIUbiElFTbnyGUiFaRE95i55JzWeDG
v7geBBmSQUAKjzvy8gdEmeIKaVct1sojTC3hW8CBVfcghJzp3kU5RoRnbvE2xOWNv9AYxhs65h/e
CVtY/2FaKhMyMnY6tJRGZKadGbGVySo0pL/ISCUX+jpGpPMQAnf2SdGKHYFU8LxJq/s/8jr0sZUN
kputpbuFagOOirRVWQoqoIG9ZRbCs5bjQ7RWvx+OMCLSXobJ0eNDCTfgBMwB5pE9gErzTu5Xcx3b
Jc9qVP0nRN4p82Ahm0oTRxOKtNGvb4ZPgpEWZOBPk1lod0bzOHynyEDnuFDQjctVGIc4zGyBs3fS
Rh7Ex9PpC+U7PAl6IUK15AmqvZQMIQy/8zlF3CuCazAVd8wlUsvB1Y2VCdZsFY/A3W5z7XEndazB
7XMIvL4N6CAXopKcHAs3ZRgQr9234xRbBTx8GV9c4GKHHNHdl0gXfrgjqGdDHYL0ZPNw4HEszvMi
gNe1vm0E/WDJluJyj7lvFpwOyjmBuFj+KY2WX5jXwl2oUTSO1ziWLFhkbEP3uQ1/zaolXyPUNWit
mln4TVcWoIswgiyE5DgRoz96hgxd8isZKJS9LP8N8uXBBVl7aWx5EPSBUQ8jRW4RuX/RAhY7olhs
A+cbDVcBFoWam1So1Hg4WLdlys5Wo9NsfmsEnLo7XuWUo2o5p2nqHNrpwS7+lLtHr3PFHL4LykEH
Zb54Sd0EgXGNCbnuP2l503y3tXgSpCts+JUNcqzuDmnEduRkh93NA3ydQ0m5fc9u3RQ9WmqNMEWR
UF79etQ+VmrQ+WqEFWeIConWYaqtR+GVHBBbcVuCvyhVHxlxWOw9lzGeQpzMrhmTtIeqcjf0M/+R
ClZSWzW38gaWHbY8H5cnSD7Tj7xp13Q6JGPMZHMd8us/BTDgm9JYF0lNSO8mOHZcjBxBSaodmaOu
rfQYZkWUaAe5zhxqIYULY5AW64s+i3gred0/jJc7lTVoTMq0Snn3XfuCvVT7ExAayezxWx9WVGjt
woJNeBUtFwXwaieCk7ny+Trs3qa/eDAtIxrLAnxJGQ+ZYIJqC8GpiQ37aHgdH69/MxktOk8+0Dmr
vLpW4hlpxCdIig2vHOl8spThSvdda8HzeIeD9ryqmscmT490r9LIGLxF3927mUU85u6jWM7s4SYE
rO5to4fTLdMJyRZLsLplQPS4Om6IQb+3e5kFUK3nkrIk2hgfPUIOxJEmMPnbISu9qvfYRAOr5EYd
uQSXUUMXXAlUITZePJNarPMh2vfhO9a+WpNg6rcrtXSaQPTBWKls6J10HJCLdcHa4YS2mCYrqprt
a+JRUe/ZgF5mbj+H1Pq3uHhmlafVopuGbyNmnSe/Sxnzk+6+V7yXfKNzs0FRfZIVRoxuPkHwhvXj
l4KhtIO0484qaIkwXWmZk45t/4wqOl5o6mbTWJBx5Q5XC9OxOlTfrZhv1y4k6Q+i/zHl0kF0+fuj
RbklMc3B4t+UNSdyeqdfx9zDmReN7cPlpwYUttW5S+qOlnjxU6/RBe24sH1ts8V/idxRX33j+O1W
5PLa0gSVKxJheqrV5KIhx8BQksfGjM1M+tBtSURRtT/WU86swlqWgeNn6K8wd7tQqAVqnxhaPPlA
YJOZgTWtGi0ziaK16uAbGOPbLM0CJdQ1paKfiUWQj10zB0XA88QP65rPOmR0SgD1EaiAc2+Wt9Fa
sGCtxwm6gPbFgnEihUXVrwTFODgsxBlmroqYVv/GuX1U+oG7fy32JpvlvIqTF1WFjXoajLI5Evkr
eRi7E8NuYPGzFWuWo1TNhpgaY4m9mrtX11oCd5acebk0FXzbS8gHFLB8quqPmSUftOwHx/ECIUJi
TsTXWuNAyFJ6MqWZ81QUY+49c/TYxyAu7RpELJDaEL+Y+jzuED02rWSmPOZ40Unr9ZmEnDlKsRL9
M8U381C96mlTfeOSdxfABYksRxxeZveWAjthMloFXKO0XhUSCJfCb0QnLrot2QmTPgbgbvq/Tbsy
jQWUEznS68zUZl6TKrIG7ibCH1/EYNn/N/UhT6rNi4CHxQByN0VekfipxcpMdzM/yWs2GII4lmmK
vo1OknVOGkbgrMeb/nVQVBNaD+lMWH/UApasjp/JZolvKEyk0UixhboIe796+7Ui13rYYRCwC6Tj
3laFiLsWYAhdgvAIvoOgrEFHC9cbbnbFsKhoEwW8RRChkMxlmwf9z7HrWURBYmHri9L+HaZUH7iv
zrB3V7sqS/5uW5csDXXyYaUTEmhaO5dSfKGsCgYpVGqwfRs0WdoTE/D2jyajYim8QxCekWkm6OxQ
C01x5VfVwvVmHgd/7jZ5LLdsQAI9QfX/CLP5OeA4k3/FLVGwJ9OeSddV6ILIQDQb+89Ir0y9eMrz
6TN1VOOKthkQ3h3g7dmZfR2q+Bb39l7nEBXsaYkPlmSutG2Ea48N++GvpGnPJ6AOBibNGrgNtwuU
EkWchz4EjIaybs8ZsotVNHoSuZ9dPtO7jvFGenU7DyfpHtIBteRk+7Ok556fT9pzur0BiIIYY7N9
dM5aWqSvEK+hqWBaJNXkZnyHY/z7L0A13TyHQBZslNFxBgFrEmS1iUo3Ds35ZiRSXe2US7TNBqCJ
TT+dESXzF2VZgiQ/OiifiJ4k3FGINiJPGiy3vtAler7WlrnOpC41DzlaJrdUCwjqH0QkRvZhU7ws
mXrBye4ejUbiWZtU/7ARwHoGB4DLA3SEtDbdj97NoxThmE7/PjSmQxbIcJTVY9p2smE5uQRKyxH6
ClF6Y+ZwBCAz0rDbu72Kfctd9lA3+OU/x3YIGbdTCSnqSxXphpVnWe4tqMMb/hZm0nj57TS6pPnH
oaK3U82T+I528YKpra5OVTP+kVBd6+69q9IjqrrlPxHGYEJstn2OTTDAXxpX+MPoolrbSSgrD3k4
rI0MBIRP4kzmhFVr0wOHNwmiRLHKOE3x0zVRDX3SnXLLRTyeoXfjn+BqBbU3vEtxGk5zVUcDpQ0e
Ql2aOfYj9aQeHUgyji3FwbxMgC40ZqyGDOnEIKxcKRDuDOSXd27TMpQfxAUYBaQiVlcN7ngn6vnU
8NBFZodcWQPMjI+bumSUxCpp6/5IsDZqQfrBv3vwZgb4oUh37DfHuJvZ+V/iMI5eFdM9CyWfhFEz
/gePE//Q16+3IfmSu+QE0poO0/yliDICoNfxdslliGQkpcMEOe/5VoRXoBySwbmi4/OtBGAdgrp9
bzBbzRie1vR0iuQL8lWOV8gnaXjwSSLcqu0xFr/fiqzlOrnoArDaRMuxWfu42Awitl+WJjsitszh
NNoeWdSNB7Wb12rxQeWeU+7GQXjbRuuBZW94I/lbWn9GNfSEfNfAuELg+N4MkFqiNmkI6Xx4g9O1
nv345R5Wq8eKSUVx5386vyP6qZrLIChm1VF/oYRMhCePSz+9ko5pBpTNJ8GsaJ27uV2wJPSltswK
rk/TQj9jN2h2xSuQxCes1uDjShI9fZq5Ho/JFIpT0d3vmZjNtsrABg8qUKp4ISlnyBguHTAsQLas
lxLLcfupKiMdxkm7zA6grER9Cul4n6mPBvhbFZ1ig5r4WWqBfQ7e3sQlbaV9+c54Nnp+tsmZvRGB
Y9EI2f+hZKasXqXUTDvvaUaZf6idZXOG9UdDXtJIbCI6oi7+cYYQ+G0PEFdHFdXBTiuN7KPDeK5C
i+EKDAnk2f3JEtEl1O5U786EhJpMqZ+/TEOz1vTkBTLOPt3FaU8P0MKkuisjKk3rYcEMs+CX0ZZI
rihW1OGpUnGLk3/fU5MphteG8+Q/3ikME8xd2zpvFzAjRkhSUQRfl39EVsInxYQ/HGTmcstXiWEt
nq59C5HQfK6y2gk307mAWjwp92avvK/PlKurKIZZiFhKNwI9NA31VbATsjpkjYoXXLpqnxRSPZ+n
ALIOKaUEigxKycI9sZD5IHWWSEDGvLl6Q3EOC2atOhDPMOSLZtt8GthIMOJCbaQS8jcRNdVifRA9
RPWyYM6jY9mRiGibij5HatSrCAKTI9hFbfuuFVIXKm6oqx+ZebItTkScVFxflN9S5ywd1RxF4FQM
6EJyGjMiwzih1V1PiXemX9sIpa881hlqC/G75iKdifJqNOQFguo+WahLSr0frffv7J3ECkj8rleV
TsnKzCMu74hlzcu3rCIH6okQMzwgwoBxfSS8PlQGNBOq5oqpQm3JMUotmThlHgaKMvTTB8xtRikW
/7wTteBIypd8yy2l15alCkFll5c5IxgcW10RvrVyVUHoZG07HfWJyXmKkonqJhXGSHwPRdPXh4Gj
AZY4ITyJirs7+YOK9t5avaTnxGRgqnKhRUDnoaRLikI4/soNcrmbd621XPoftGE+rPsQPi0eGZe+
t3IXqaX5Nlr3dDC2rd3t81OU7Ce6LlC217Qc/FHk5KGVJTmilqEdB45LfRarHhuDl4b0lD0ukNu9
9RcEqIoXYCkmU4TnlsRLBFr/Cek0Yz3B/aN2Jo6/dKn8Fvy19DyTmzsyyCohnZaFpHwdSnF/wOTK
R8H9Fp9Tmd4+setP42zWsO6UXIMEdZv1Hgm+rV+OHrFsupgQ18Phwrz1xyl8bmmUk4m/5mTKcPuq
qumC22MeVv6CuSyQRafwQlJRA3QrI8aYXKNiaLGVCgbB5TwR+OIbcv32HyIPWswvRtM7MWsnS7hb
lryYdNGUHN/hMmFYm6jxDCEesqzIRxzrgFEj/xG7hy1j1fnu0QeZZr7XINJFIEOedmiPvWCeN1s6
DNfykYvEJDFBoBkxfIQPCFpSlkFh9xGs6QDq1hXNCpdJyRgBK5AXNFTYf3HS45hf+5LE3sT2r3HJ
ZnPBS37/T6z/wlRTGE4gZJi8B4TqP7m1ye/sdNcufnwV7dbersContYmPUiulB/SkDaKJcSYDyR8
RP9YlNtxQ/eQmCVyMdJFQzOkdDOgoXQB0ra6hJHJlfGxuXx16MBzvV/AwSR3tn/xVNyJAvwJoTwF
e0S9u2fqg4WVTqu6Ut2VvtvHPa5gMBVLdQuQEtzybqF785N32GE4Z+KaBKAQBMWQ/tuGLjxbEC/w
1QsudA23XWYq5MFriUjk3/3yBdpE4f4koArrw9ZXh/PK8osqygNI3TvUBmMpGZWmO+AqKHBu/n8Z
KRG4sV1vj2LUH49Lp0AXbkSz+g1xEAfQaylDIQLKelJaLzEMGXRGWRao3Nb9O1mdX233RrztWwCJ
Nq6ML7/mFOmmd3AGpHBQB4Xphwhmc4BKewFcYWH0c3pI5esueUPZxFMl9RDaw9hoqwsJQwhmOOJb
tgKq1rI1/R9gFHIJpddDvDmbElu1D6dafvxP5DLsxIR/BZ5rbg9QaIM3AIPAzv6wwH1lEdvKdsfu
0IBVLlwQFuu6s/DFOo1z7QDqVX3oDN9dc/vtQYA/2h2M4/2B4p1HWgSZncB4f9LGIw3H0IiBBRFK
x5752F/YnPqvyN7c6ZlwVK2ZhCRbunbhgUBHXrUMz7guYdImgI1APXH4CE6XRhD7Q1XGwykDEo4O
vhsh5mbNKoHgjhJeOxDJW1YY13+tT+vRIE5NdgmyzLJMtNnIAVlhWMvkbYZvs5N08ugnvTuboClT
CxoevttQLCn9/hWS4XOuO6uVt0nRS4sY6l8ChWPwDkM9K3mq1tJeQPXHw5hfN95aQxZScDBRT19n
wF34eNGppRKqG67u7etzQmT7HeS8l6ZIyOEYyen4EymrAaigTmAiXNTIeuZibVnkL6noRSAhwghV
JvnJKIjykKQpCz4nqxxr+aPR6qPhfGOefoDU5YA4bAq86MYWC6Iqmro+iNy3UF/EtzdJV0WOjjF+
exsiWN5CaAhd5A8vnn6j7zqSm4PASUrabS+nd3krr7+bNk68vNvoNrPNgFNHBfNb4IGhi9Tiy1Y4
N6C34vNaCigou44oq8pRdJL4DNmR7KPGt2vm/zaO/qc2cIYVJAD5gxRU6LwSfpUCehwnvY/u0Adu
YIW2Z/+6WABkKjBa10oXnEnWqxCwrpGuHMjcjb/kNvbXTvEKzOBjAAknA6WL18cEd5AvZjo0CP7T
uTYsP4q5tC8TJPNcmvxdhOfKYm3dz3vedF3p07GtlUSCZo+DMjaDX8IRt9u+2eGzaomLV7IrxFi3
ckuCanPsmLnAWAYXYImPFo0EAR+yURB28ScG7d3/0SfzNuRUOZ9i7WhKR68EMStk+yWllXOu5DkC
cHSg1tP0OOkg43ZsrL0MPlQf6e28iZEPKSKoQ1qt3m1ySDENENUrSyTdqlrNbP3qzPK9zbxhd1lL
oBifpxrby0Z3VQJoYyJm2aAK93kX82pyxfYD1KBQyI+dNOFqddKAoYbJb5qK62hYrrrcBogEFAOb
VKwBAXsr6XkB1X/33AsNoYoHZxbxUqUJp07TmLLRCXvhtzx8np/PboTAaqT0zWjInlWe0/2Izk+A
P3HZE+L33BJ34fs41rd2JGofIHngNnyeaVXg439Keny22KCkhjDvWVbbAjsYWD4FiYAoWhi51b7R
OTm36zUCzIerV7CUip45CoQFxvK+cQuWsNgHTPOGRN476Oe5pOU8VaZt93Kfr/C4GY+svfRacus7
3900MYG+QouoJtesNfB2Robzd6r0cBfvUeCwv1U92GQqoDSgWkN/49VuqDy+kX/jMYHAQiokNreX
Gc2ql9WXuFBgWJMk6LcLTByOD1bNRtzmi0veobKtsme5Ht2OlKmJJ49W8tKoOOlXCHW5IPpQRZ07
npJ3w82DQci5n4cIozTYZ9TOdom9gY1GzLe4cjbCrdlFDqANZ8xTIGZ+L1iah7T60CarSypzcHCL
dlMqE9gA4QuUWJpHHb7Hmov/tW/NKfPPBYE4wrCFu2zsMzEtOtv+uWguKHFdy+o4mIpiSVn1ibry
tCpEZSsLpwvWnZnBY5LkhP6QyN9KnsDAYXezyNttW6miu+RpbYaD05ktgNI7tK6R/DJnP4bUwOSZ
753znBJEKQrPKyCuVvUTxIepTI8JFKgR5hgsZRDNVikqeg0KG5sKeeiTjTcewTWy490wih+9F++H
6Mndm+dfztCDETuO62L4E3W7wIMYP22wYA3J05hnIYJcA3t3c2wl4mgfQlfGGlPAD3kOFIND9FcA
EN47+rTCa5QxAZ93/MzQai0623u8wpSCybe9RxjCqGuBRONNB7bP70gS8dgT0xlC1wQ42ntTHZbw
xNoGlYUT9rnjYr8jtMhq1CQn2BBz6csDX4N5rqPtocXgt+aYevqyzZhD1AXu3fVEuaIUXIJqvh0l
VLWfH3pNRHV6ET02LrwQECMtope0ZiqrjxI85SsuvWzhSNuTCw/g3l9E/TIU7+fqM4eNp6xFX++B
cyqoEbj+Pl5UgzKgcrWT5IopduaBRa0QJNH3EfOUVXcRzG8DMu1y6g5XmxvmD9w24WTY59oaqn8M
SAkO98cbqRca+w0m1heiSwkydnr//jQZppfGV9+NBCIsKBq+iV6kl3Z4SzVhqMUOhH9wDaI7R4Hf
SQ6WJr1XakcvRqnT8b+dcXPCO1sBkR797dgtgQvgUtqzegp30h+4qwathczj4XFJvbhDzv/GKhve
PGH1lqYDMmg/vTH+TiLP+0Jk7geDVlMfD1J48ONQ3LfvojnNoNuSSDwpoBWAzU0fPUF5yCULD7t9
t3jla3A+TrEcKbMYYh9rGmKsnw3bTJFlgViwU7kbFhq76c9XT4+2qdwuvygxR3z1qZVmbcquZ+V9
kCXUgHSx3HddLWX18aLof2D2nn8g3hfu9OLp5ETStvv8nOu63pnb7QrNrjer0U7RYAibRJqlTAy1
K86yJKHCuHtq2+/1C+eTAW+xWiuhw9VvBX6DtSCHgqPRNYVw8DzQJvFxIQDQt8V6JklPv6wRoSre
Vfg+NFcPlka8l3jCxvm1qzI+WA2z7XpjBbVki83HDiNi0T1fT1J1QK8NJ6F+xXRFS7rWDxAU3YG7
x3nOjLA6nu0J0CWYoP86yakB5/KCCkgFmfXufNysEvNyH3R4rdWQMmIUbAOXGdq40x2fMQ6Iw7VO
HALOR3Hk1iUPv6yuy2vYepGbzvWlnKLna+cg3WdIHWm/CouEuydZkFzMb6pciN8MFYhEh267levt
np6g5CaNsA1eeBzjXXICVePd3vI5Ys5ut53EXsRa+MzRV+GORR6aiea/uSQh03veRE8M1H8wVZqP
IOY6rltlkmQp6niFIx6qQOhClKvniF+HU3YWZAz3IyI9D5w9iidNZ8TXDnKp0YOetQOzDRXghMbS
EC33xvWGpsVx4txntoIKccBM2DJvW4NddKiTAow5g3b9WLGAVIe/vXKKmBQ5ORv8c8lT2VjKbJO/
qQIkygeh4z1gLmFWBPKPJZZVCxuyhLw/yTV2FK9JgPd3pCriT/MevHVU7xiqpMqp+iNU+ruEdNjK
OHgIj2uX0GUg7aZQpzoFzQnlz9v/iptcU+xi5znCe0cNDxel9pJiWpZiRhXASruEu6ZzFot5K3am
8p8LqL+I40wM7vnPLLXo/JmLH3vzBDiwXajCwL8pwc7HUU255yfHtdmg7PLqI2bpzngu0pqL/FDZ
XRxXe85vXEv+6MIylLC/1BCVxUNUqiD0FCz9Py7YGL1Zzo1XvnbMPkhMDvozjAPXQsLE6hdngdkC
bXteg8sSsCW8CqiihhpbqLsdZ2kOn1sHQpUcbZTrrETa3F0ppvRKBjUaPFaXFIOisnZxykG5Axpw
fkTW1t67qA9TW/gsk6bRO9sFLjGfmKsZIzYPjdLzDT9hhpg9Pb5Mq3s5n0ECaVSOcRvKyfF93tNA
uj91sDbcy1E6v/egS+h00iVy2bFYqVaWA45RuApjOvlc3/DELWRW0yLW5Fbh/8h++sdq9YawWIzA
Hp/K772S86IMgUUnfpSsLGB2PNih9dedF8p+/eTrfTT7rbsZztTDkzkmAXgWMr34umAKjfqbh4mW
tocI6Umb7PERQOZI+nWFkwoLQIX+aelr2knm4X5glsYEAiIe9fGlqGp3e82quzuqKbQseuCzwwRj
AuxlBA2zNZSiLnhhvJDS6Emzxji73RLfeTnc7Qkg+eQ+Yw4HHpla7cYxIXVbUxtqgu3TsDOfetRu
OCtqFS3rQa7IZNRliccjcYNp3CYbNTnFsIuNOHEddiopW7pSNnUej7P4HHQY2dBCJFUedv89k0p6
7WCkBLqT4qE9WztLFyIOHX9pg7bi9wuKB8PimtSPV/xhqGW6JAat//O0Jjry7xMvsZuZBqIfwK0k
P/hYHPthcIhPgqzXR1jcobvWZQoUDwzXAMphgqrQ5/XcTfrGYr8Mg6kRvTk9FYvTYAroA03jWzcQ
PWJmHH0BbXJqB/nq8dTMiz/sTZM1xxHz4IkgAx6FxTfpUH3cgvx/AzNn5T1crSl+rIUxcIFJLW1R
C3zpAMR7AQ2M8qX1iAF8fkfl4EcEPiqu81m0+TVzzGJa8Aq4lpSUhYBr8soTKKxYyGKSN2ZsLZoi
sqrx8VEpN9KuY8TjN9MRMeje6bwlP8Obop2hQrZidiCB53FY/4e3BGecX+SNDdqxfV887MoOMjvH
5ImjVq0aqm7RHJm7Du+AVEGP166SvNL1PLO/veHPJh5V9R3Jxe56L84SFI/Tj/M3LJqb94OMThZp
sGtYD0rGeFiEukiKHNRazCHfLaaAQJ6EvBkqHrOq9danIsBWfFCd73p0n1e29h3SImKclXk5qbg7
PZHCYKuXDrkZZ+5htqA8yAKMKNgCV/Ye5jfk+Z8vBfX3xu94D5KR0Jt2te9rjJ1sVncgvDozS3Lf
nVdObyVpzTF3FBCPwjmyBpvULek/SIp3IhWNV3wvtjH+Myb8X8xCsqiDjSM7LjVv9Kf67ch8enkr
ZL70xnjRk+5Iu6tPFIucRQobXrxD0FQnJObrIFwAGMOpOc0dt2+1RZL3D9EPC/WNupUVMSWyKftJ
PoIYl+tS/7UaGGE601YhVy0u2KhnwNcNacdUP2H9pPwEd//SNmXz5Rwcs74NBFHlEb+fIiXQlyOF
w4ErReCUemQn6sPp9c67fWcpSPLHib1D39mENgOuibLccASB/N+/DvkPI4DHhD3xXvq2xbFnS7F8
KyMiYExBhJn7camHJDto48MyKCEAkI9Z5OdbZbO/LV1xDEFi7ZeqH+AS6UnkgPpyc/qTGWqfb8+2
huIr0ZarLb50PnmwtNmrLlfqIHjPwRivsQ+Wey5qbhLrkj3Yl1U1rlDgzQa46dY3hkTcQ58Wu41R
GGFHO6shucA+QKWYSVPdtE26oYE/8qolxgIoJ0CmqA0aPA4q22pOHmAGOmtyZZLqyC4tvaTOMuh8
MR/aZxqGznZRCtTQZKNcJ4SDTTzQxHn6Hgbl2hB5XZ+TWpR8uDtun4Lj5clfmXjhs2AHVC7+nU1Y
y5JKvTkWfIc/DQOACcfYwaihIPEG21MxvD3NPrxWy+L5ryB8uew2PP52Kh/P/np4EXz/2hvfSwKZ
TCzGO1AfT7/6gc9fLM+a1lbSE74K5XB5Y1pXY2zxSi5nZtkY4heoWE6uYmPCTSFpx32yOxmG2EHw
WGv77fUX85UVE1ACfexM4khAjWL4LZ7m4+hcD1/NHC+fM30OKl2JJULNW9C5hqpTwM/T1rYw7K7H
/MPNx+uvrWDTKIuAO6jK0QIMEueutTvknfU0xD5oLL0eFWC2wQNTRJNqLTHdPudVr2YnXQmcLuiZ
rtCoue3MGfjfOuVlnszfKjOpz7c+wCD0+CuAGGbTkeVKI8jwPACiVpzjhT1ZEVbfrK/XMB/qr15z
s3XbA8JpGLv02grLox/erLItz7C39uLr/ZAKNRYCIvw3YpOB7uMKPk27fndZZkljDdQiK1EnjAmf
TwA5f4yOU1P1iitCrgoFDcFqtwnFRf3M390E9kHoY6uxiP9SVLyuKcwNMJJviWEDobNvElW9GcOF
WgrStQwy6taU7hETpDMwXXiKc5Esu8Slb6XwGzDA+5bMvARdUb6ved8kJ68d7aUZrQ2Siq1FdxbK
TdmNIaRhBDSXVjzTy8u0UZrnqs+CbXMbdJqaSbu2LKSdYWsaGc+zZPlmulSSlc/csUTSF53McN+E
W2E/pgORmuFS7brv+Mb+q28wvAmq0Njq73BILXQolu9FhcsIUq1HtqgPsFwfVt0IVcXx/IUoM4kR
sZmK2UjBLELDN7cUFSdw18/hWa7/7CTH5rtjp/iD2lcbpY4XvteKv/6IBMW+yxQQPQuInBA7WOcC
1ToVcHU+bVUucHLdIYV5o8akGifXYchdXlGCghtjARF5p8HF8YoPypfysvKuD5/cUY2XZRrtS6oo
jn7Z1kmad8ihOM0ZuDLqR3Bb1sDIFEfSb82Qxng0MX21rSP0EAYu/DjsWWmSZyP+kvuE/A0gXofp
3449i12tm/X5p7hbEs+uxRmETH2OofVoYdPNi97hEg23l9I+x8KuWF20iSrzbJqQP/9gngvHSnZq
2U0BF/9H5p+a5I5fWjf9/5SXMpV52pgBQamQBP/ATBJX1/aoLLvCsHHroK+3jNnfDIPzleghZhRn
DOb6OudPVPLY/DvfYF4QAChsGc1d8ZwuJpVnawtAc/+YGbs8TV89kSnpv54BkjKJ1PZ5otwBU+TK
FsvV0obl+djSyTZDupGumaiO0L8X6gUMneEsHS+3SWYFdU6ytNT/nOxYb8MC16IJUVu2Xu/ocsQ2
M5l094s/246IvdbzLveZCod792nvs0EyYh4s5gKYvGvkXABcvwzmI5YwIkoP8u41EHSHa4gbDWFI
ocg/gU34QlHroC2OdCDFgTTYaP146TBJi0GsrQCJQsiFumgGHumyyaGhgDgRh2gpZgXFNY+cdSPe
DDTrT/O3CS1i3Nefkp2gs8RboHaYWpMx9M7Q8JoRwTYX5+5I4QWb151LQtdi/ocrS5NOeYW0LAvS
QjbOM1bSHiVLihQRMwfaT7lyC/D4U1ncGziS6ep6xfgloINb862cAI0HOhuvsGc4qZX0OgGk6wx8
CrRnsNluKb8hNI0BsjYPNzYUXt6p4Lrufa+3ZYKwF+zKRj0fw/qicjrkdMNUr3FPopH/pxuYcKKN
BhNe6Wz/BgYdmcvcLkDHzJRP7BZo7MubEw8icfT5Oi+P8/MjjUspPnYD9L8diMJxZy9l0DoKeI07
RcrmXEC8VaewGmdJZvRr6UTp6zsGS4MWx1TFY0XD4fAtmSudjzlpLAhZgChPgf8RkdqFjVJyY3BS
g9uzQkN56kIVbRqav9zruy9/L6b/Oz9EHV+pzNBir7/xYn9FUL0RD8WKQoCvcA1bJ2FAe4N5cQPM
oaMB9qj4qjhFMJ/UQSsx/lLp31c4mNT+2MaiCOR7alXvkARdgBDLEjG64ggmd7nryhaxNRElXjxB
XpmO5TXBqo4igC/R7Ds2Di9JrtdJCORygPt6fVroMV1QUHRTlpViDk5mJJirBj8YPb4DdbUvnvik
OhcPjT/tRj8+gWr1GXqHuPmymzr1bCvQmyTcfHkGsPf+0PsmIQ+6DZUZbQAmr+ufl390Q7+7PiSM
8wS05Utg3dTrCd1mf2Yu/G0WNc89MQC8VWwW/ZhjOBVERTe6nbQpmocPMAa3fYu7bz4YhfgYATBl
LCovtbOTHtWX2WS+ugY9YwYzGhKLIYdSn1LpWYEWyLR2Qeu+hMVC8/a1dGDhazdnC89dJIdvx2Pv
YUFcDSVxV6A1LcWbrvbiNPgzmEwY4WIvEtSQqz4cT9GPQ3S6A47wUkMoxqOjlZaFhQnKlFsjTZWw
Wn3dHYpqvcHu3MBcSVLxjna8N+PDw/PfmnZsTQVxeDpswcC3hCE82Qt+hv362geSot2GoJw7TdLl
/F/2cy+VJRz0wanVbzEu1SJpqeWe5cEITpuSgbyk2RFJshmLhJRaS30UNGNtV26z7fVoYr2/XLJt
V+WcAYPYBnX31rlANFlPk7f/XXnYIXNv6rA9ryFjQYCpDdBG9bPI78GHilSfujRo9B5X5kZqjpfJ
tyBG3CW23NJAtMVhKdCuvIBum8YP7ee76WmqZrmV9LlxoAMYFF7O43/VIXhtWxuH/xPQsNEr/tg/
unt3dSQglZ94r5623hXU1JgAsz60qJkCMu5jWgySi/enUdbPR8jzA6tux3Yrj+UsoxwZXvDcois0
D9wK/dbhI0gmToCA2UsP2D9bAN//UZYibEpnK+kOx0UyXz8AnSjb1ldUMOhvl/pHof6tjh471jhV
GuIwjpIS26myY/MXTd3oebQeBX1WWmdKkGgAVSKRz3jYqcQ2PpWJUx/P37F1DUAwzBUBNVemnSKG
MRJGvHAntlKynaf5lVCub+avaFKkj4l6u4fhhATUQKmdtRQHv6MPXSmr3orhurRWdR4yz01AooI+
uKkhOidLp7J/56bCPrDYdquowpoTsolpYs19C9HMYhC+XQDmcJsUaTQ4kjqcAdJH9QueeREYU4sA
SC9dqTjdJYfs++HD8f17e71RB9oq0nQYM4dAD6BVnsHJOdbti/4uYEcI6mioWLQtNH/bj+v2Pgmi
dKeLqU2kA1hRdB9233XCitTNh9PzqAgnjEyfFokFJEMuj5KyMqaEsxjEQzOWbSpny5Aydw4865ne
Uk0YOLI4y5IQgc+Lvi37Ciy4AgHcmOiFsMyY+o9JJx9TDh6TOsUz53WeTF+/E7I7MVAx8wry+MpX
7QtF5e2idzWH07NwGXYt1oP/fcGJWua9Objxb2NRIC3gFRQj6TwyFsT42VQQymXyY02hpdZEEAuM
Tn2BkSKfTIsUnbCQT+ZQ7ljfMi8++wekVMiGbBWYRiOIiRJ+Bmmpyajqjqe4ZSe8EonKF0HiRi6L
6qOzXYM51UxWLOyQ+UNGdRyG9EFwhnpLEIZd3kPepl9Z1PjK97yZ2YypGLBLhXfdshqG6TlOhcnO
l92bCDjHt2cCcLTVX7adUPOUn9a5gFfUgOn1a0W7Y9lORVE3msQ21roF4T4nFl6R68LkgFuBlxRj
h4MqAXdSyKb/OQd/0O7Ma+MDgIBt4NHln3k+n1whbhEQUwEJItayChAolKznlsG2HYzQyhr2uKIN
KEPYf2wHdWLLDDQb0Fv7EaF7MCQJTQPw6sbBvOaWPHUnkjlyAgs4iN+gKH31qJ5uk4bV80uNiU+D
DTGwU6AE7DSV1CWxqD4V5kXyVwPkQERor48MAbEwRC6o4dr0R65T05wRiuEZ1ul7EsjjITqpcu1b
qhWhQXFLUG1s59ZKZuKjANEJejEc7ATQ5PF+WrdWgsEnUy+TF3ssrh1OSO+QJml6HqEPepNeTwYZ
7XvjPjYXIZeAkKeQMudfJp9DLBu0zLC5ogumPig9oHkPHXxVuEwIvVBQSdSja7L94JZvn4cf2Jvs
sTWdzHHEFqff1JEJtVv97y3ErTug3Md2rO8sDkcaH6GIfbjzJJGz5JJtD+MQQqTovlvC3/VFuMXT
1YjLQmuhRIWp1ayjzGU+4npXqxQ/T1ysK9I3QrXkMSTeCRes8nAhd7Er0VYjnlNDD3ViKKYfs6nM
qM6YLNB5o/PSKG5/Qn2vDifjd1omrd70m/1InEjjtBfAyFD0V2aLikQ76afhVmZX/xi9R9JlZZA4
UsCkw+I3KblnuJW2C1ed0xjSoPSSbyIhLfhdZWnSNDTg9jVTyvpCIpxwb8O+42WVo4/Sd8Ohpo0D
93hGTtyJr6d31dv7t5oNse9F+LtDwqqEEHtJd5o75KClpTtvgXj+J9WGIg4q5teABA7XVAbc6wk5
9cdaW+A1W3m177F5l3eG2ro4hRqegYAbtoWpLMBYL5xnNHSKCkKWOaeq+HStfzUvHO++KfIxccNO
5E4hMlbyH7PzZwUXEgmfLRua8NKUWpp5RlwaB0qkSj77cUAFoN8ijFfDkKwdKgHFzlqQeEQlqvtu
H8XuixlBTKuUNXHJ99zWdahdLvlDW4fSZV2PTI1oTpaRfK+M4herbdrAC6KM2bwkU8Fk1f1v5PBd
e6OK5IZ73Y/vp5nE/hwD2weamJ1UhK6Y2qabLCqVs5TE2u9HrUXBqmtg+N0HWzh4KGKT4zFft9WO
IHbIFC9d+UWYa7wmGsAH/OtzwDz4zMDcNsIDMO9dI1l5FJs0HadYoraE1oGLKaZlCn7VHAqS6Lzb
YGiEaWKr+jdZ/1bFc4wLOC5dP9H+tbLU6JpZfWZGqEgOPaTFxg0Xh82SMMvicO1t0zktqzEPSiLt
GVdhiLkUrNldTITrDiZ13LliO//CYqzrwnoB1eZtQehG+fwOrRr3rTbEYYZEGqx4WRN13e/GdUIf
KB0EybtiKFCDn3HiNmH+p55cNiJtj/a9zJL7ceLhhWSaIJ+pWbroj5ZH7HLrR+MC2Gvdks7KteKV
Yu4PujYIOK0GBwlbWa/DWOHBTTWPl1I8WbW/ZXzKGBkD6OPT/LHbVPgVYyHbCTCbY8yIO7UuioxS
uq3zaZ4uJMqJrpYwf4vRWhzJ2MnVgxoZa+aYVuZP3Dw06dRhJiYg9Fr3Y4/7rzvOqo6jTxX2oIXO
A+EDqffWFv5lOGITCWx7y/IumDRekFgbqMxMYCAiY+RGbFwlTah/X3AYYoZU/YJhLHTnZcsdmspp
bfxz6fwPWCPyXVTrlA1J1mJsaITIZc9VXt2nGaxx3BIlrpHB5Rfgr3Ozogfk21/Jqmcy2SPXD+ct
cQRv3l8zWrFcE5hxk1q5tZMD6B/UZBy+uvurr5gRHsUC1YORKjeicxJrp3ieCt9LUiuM0tiA4TKA
4Km+Oi+ikZaqxf3Tvf1C8D3O88MSyqauIbSlF7jYisgnwz1kivPePpnNso1SLtT1J2+6mfrQ/Vn3
erCrWJvgczJ+++SJUkKiYDXhkUBJ1VZDAqsUPYRtmjsN07XcDUnyPe5lRLepiXvaRzrzW1mErpn1
mexWRAkIvsYYemmDttRN0KQA23vLZ6Wh/v/HODB8Q8uF4gEdhTXBgi9WXjamV6+jipBnxwS95ZaQ
PNege47HXEv7aVhQ1/OAdHPZFx/BRjl3w5r6wUeZkUTAQxbYr4bVy2x2LqDenYh2V8VeSLvc1eCS
uDimiI2wI+zhIg/rC7SUaqAHz8LLTqoEAJsdd4SxDMUWK3p9PJX8gglGEgaQTBWEQBlah1LFJP6d
NpqMV2ZOiBDLBXtaLVXGNqcXzXS9NI2JKgoNNrZpyP1yPx/x6qVhutUH8tqgOIJ8mMpltil4/eXS
71NG4z42/GTkBVRevDCNIPwMDNvZ5LTf6+lWCoAgJQCXlCZX8ax5kyLXKSwMtoOC3vwJ8YGLN9ht
HLy3SqcXqew8zOmECrnMRADGHiywBYBr6JAPpXA2yyOXg1YFQdFtz2pn5nkz3RxXiNC1nxIkOYS+
DdisP/UQCW7qE3ih9ZLNN7QkrlnMDmZ5/bWPhZ9mNyXVDZ33TmKjNTR1juRlftMz2HY4VRYMgHTF
v2Rjmd3L40rbUINk73hwiHZxQ3DbtjmvmTmU7UlfsrBo8KP7iXd+Fx1PnybUD2FP2wbkFLkVOVss
FDRc3jZ+2gDu9MszO1TvsXCY5vyoHoNIFv1vj2mfiPDyAdElRaoNaVXc5LOgOtLtxlONCs3Ay9Ov
3de4Fe3fSxcLg2YwCCFVSNpKePFQ9bv3R5/XVhdPUmm6BG3Pt+NxHqSqKmfpCp3xsXKPWi6GUzrn
UKgAX8U6UCoHUWekSd2B/A16wsz+/2qWBDwDaMxvl4DTplpTWkOtnEzUHQ/TKAOLQzfXRyt+qf2W
/ilbwJ+4mG8u1995+QrPCnDSXmStHDDTt1g9t99/mdoEz9C38RqXB9Gyl54IhKCXm2AsCXjS3WnW
jqLSQxJw7KFaU/3hJRYAsHCsLI44vzyszkZ3eAvLcrWL3d6TS8nuaQ7hUbEYehc0uQneoCRtnclh
HvHFH/7rtMn0/Au3a7zaWE6lf20AJLpDrXQGgNvaS+63Ae1HshDMQtaF/1+DB6AsdFreNOh44X9K
LZQ/T9uMcZXcFc2TZ5i4+GXx39fOK2qYcfIuKZNVJfD6z1DAlFE8qRoSjtIEKJGRHkBTbsaq1o9o
ZwAseGWFZyrTUeld0uRQ/wvcCNH841n2zFW1LECg2Et9ArMeJIq64Vqj//it3vQcoFRnfQJFmASt
vQ3Cu5uCUo+wVWbEMuBqLKY92sP03WGZgOTTejowhSWcQiPmEaN09So5hiMJkMWLp0NW85J1jkVw
oErs8oDP6YohRye0kEreJQE2SxtsHSN+1y05JIb2JdukxDYP7IPs3k2KdIT20KJim0p6fO//BgUj
SruhqEsejQCTptjlFZ78peDM/BwWUI/7Ct0kxNg1DE7jlDj/BQ1qiDOpIX5fsxa6b6kn98q9TwXT
uNYlApmgnDWnk7LQdhLzVm0ssDZRmaL5ghBtRthyI19ius+9jntj46+6W5kcap7lTb2kaA6XmoDM
YDdo9v8uu95zo1+l3cdyykCCQGOOtEaMg6blsZMSAIUV/Evi3zC2YpkzncvQ7uRKabTL/pw7ZIy8
AHaPxFLpkZNjIcRw6cgThDPZMtQnhIHo7nHvLzMStjOxSItX5LfOl9edANi2UFCVKzopWs63Xltw
Dh5T4Adryrwd8bZEpm9QM0APsDReuVqJ6e1bm+E1Y8N0Mc9DchPe0SUoZx2tIyUFB6+N98yOaOeS
oDIZ6MTj2ufN6+2Rb9kly6kG8AoUyqL2LyQ64PBkvwE3/M/JStE4FK6oza1CPX4Cr0+fWBwiuf28
Y6FhGHFlXubKiv822t6mAlMv8fWvwYvVV9DDU/BtfP0rcNL5KeiyrKUZmhj6sJXLOOHNkQq89aOn
OJWNnsHj0yZt26eo82Ap3pOQlmCkNV2W2w41FpG9wKG0keZGFKY3DlilQz/STWTiW0oBoUcVuYXp
xHtlZsJGmyZNcikDy/fc+73gNx+pRb3qc0oqwbuEbGwiGr7Bu/nr2CF4en2keiqmeA/P6fgtzTxF
IrRECshPJ9upZh6te428387KeekHCiFIAw7qrSwzniE1F8JihlGnHeQ1oC2CIUnkyDkEd+swmJ77
/pVsZLzDIuLs0icajRbHKnEM76x4VuzO9bK3afWhrd+RRXiwvLcmoE8La0upbaBMfdtUtDkw17Rf
KMTvEvLmamkvD48CelyglHpDak2+KdtGt/TfQZy6/ehMFJ4y0Tp9eSH0BJO1Ak6epfsuAun5jmMS
29m31xMXSorqD2CMG4/DAbERbfr0IWmaSi7nvO/WThOEyRDrZPdt3uYpj+lY1jcuAEeycZI6/mPl
wyOnyVHyQ0NQ0SluksFNJJt6DUBBjDUyyV/+8yHgv2rlRBIqJpsHhaFMgnEk1nOvgOTAsWaph54N
i0owiHXyF9+bIYvC8BuS0TZ5rLabRbh8hGYjT5Oa33Tar9kSA5CpB7zTl6D8NYGSKViQATU357/F
9QWljX344sf6AOuieZ3AfsT938CvW6yt6haB9OfzVWzxRZ+OsabN1R9WmLA0zcZCTOjITUywVT2c
yj8uNVut1usUZEQ25nzSaFJnl7QOsu2ts9ikS1FEYSJCe3YIGstXyfAABjzQpGbUBScD/wSSPZ6Z
R6LIwjCrU+pxNreddFxGg0p8yK1nnQ/cWp+oszn3SOkaxWOz9TB8FweOOJcAt0j879u75owIa5/j
3eZKmr7N8NE66M/Nat0UV9PBz9dPyYvWZCpAXGNQ8uUZ4PlsIAwV2AqSBE82MOki5S6dlQhrln0a
3JkvkCiQ9z2ZBXALMbZ0AUFK2rKnSq5GowkeuCurAwc1/jiaeoyTxVHKKDiPGCFYBzLhA4ht0P9o
xqOL7W9nw2sxmI3pvy7kxexhXSM0CudIrZzWIXirfKMp2q6uMldvsC1HVy8HLVVCSSpaBsDcztgP
PxqsUjg6Fw13y6jaZzjAK7ZXkxWWHn79ola8yvFuYrMWPel44pF09DulgJolgeOmrhoJRRaaZp6Z
PubuKOZZrVNtdMRp9tZ4BRFD5No+5KkEHlFkXdm5CVjtP1Dbat+ml+nHB6vFL68j/CxEhioVeGmZ
z/s98u2qDDW/9aAHm6u/U28EresNEGmYrU3Jq7dj23RYga6IpHv5S0e8VdC8/Qrp8REREDuEwRfS
u8RKZK6u+GVSBaj59+869O3oRVGfSOs1F9hYJo03IyQtEMKQlNzDEXl2lmOCyF+dLwEefzKhgEyr
HgNJkqoyhkT8FBlr88WbIOErMy6PUnQUPAhuHc9eG/2CHJTzjIw5tqo0EkZN1gHkXwJE3+xD/RuS
SE/yw/H9ZYuN2LsM6ttfx87pFbKpXP5oQfF6tm0kxt6grX2kQSps01wp6Nxw5Stg6ov1VS3lp6kI
GCBPrIgrsHoVooGoB+uEQ1dqgOdlt64V1lYVUO65N34Qt6u9jv6cntYxr0XtJf9WCwYyOwsn0JfW
wim32LB8NVVF3kQgncvAECAeMcKvPAn874+95U+5a8VBs4T+hbN34C0kmAJ4sPgFi1GqOyK2Lkxm
gavQuxtbjBO0oiVEc0BPUecdKEtlaQKfql1aU/3tyYRUWXC64+sP/XU5GvKbbnSC8NDk5B5EpJxX
FP+8r6W2AaBVNWkSzoHDas5L0iRhU7vGbbMLh7uFi2Qp3Z+sYl4VltAQX0dOkAAR9o0eYTFX3edx
dO33aIso1zGxFsEcNaW3c/3BbyxB/p6qKWHaDmArDdcttkr5eil9k0k40R/N+IfmjzRPxTK9hA7x
I1jVgAYBaGJtjtbkYc0lNsTFI0dTxHR1cIgFfYnUPWdz2Z2X3hrHTxVIWgYOJmcyNU+Qhqxzhbk+
IeuKxp6yksn4bLDIHSKbnQrmtbcI5VtDTr7Y5RTPJxJLjK4IA71Oac+muUWuR9rKDPEopaTe/x2I
EfQzuwRoi9a/46PQGvFo80dWi/NGn+Vio7P+l2RqUrd+L5SWTPVLHGCxcSJZcMvqKY/GqeZVx99U
d8Sg2D28p/Ns9liB78DeUqrIjJThxqRCVOEbm7wHm6c3UwNlOMH9ZP0jduRdc1uKnudpPMmi7DQF
8Xl0rWqWR1Dksb96YmKo0WGKVaFgNRxy7kDajbYYnlvEqC0PHsAsvLMAfY7GS7TvXgqnmLTaI5PL
iHrKwzWCvJOmjH87skSq2gSx3njnF2/or8hU41fNTCnOacT6R14SijeJC+vRBH1EHn4cW5/F/sYC
3Mz2sPajy5aN1/+OQ2wlLLxU9YXxPFSef6JfLRYubPR8Td9No3okYBNLxIq0BOxwoWem98nga308
d8+/nPZFvLP9/zTQKFigKLItjp/PA/jsDmeUr8uowCuhY+sK4F4v7xG2qlf0ZB/KC5uUDuwUTkyT
7AbSrOdcgK7AfcnK+H9DUthappIGMcQKorz3pMDC7Uttsv2yQAMEJ33U9VmVf6WqeO4VhMuaBent
DcbljTWb9wWI1TVs+8/OAEUBTswrXTiJ9iEnheok1Jsot6GuJV1hdGPqHxk9V/EpEE+8E8Yidp9E
K3Ge6rNo/8darijCVcmmfzuUl+LU1afznHOCcnInBU/4Zm7wTaLWBAIdzDjdaB2baq5TJmjdIXbI
RH3VV/F/Q+2wJkLGI6qv+s4Yj0GyRC+e4Plvnw17tERP7nSGniVtSZCbxFmJ628MeeFMxBfte2EE
xnGIky10SJW4UTeyTLCYzb7FHxAAGtC421P3dHZKdrzqaE2lyx+B2RmQ2X3d7KlfESqTB8IML+i8
7nN9D1woTL0lgtgn9NTiFPlrGwhRVcuBdlvt8HmnulDsSy46xWDqs51wqzYmm0RR1M5zyFYYuBUJ
8hL+LSVtnVkVNaZvs1XD9jX9AM2efzG110knzYYQPnZdAd4LeVUNx2j2hBa9eiK2tTLXMoZHLjKg
2h2dC6trEGOGWg23c5z6kH3DTs6Y9yUoyeTEwVwKegGsuoJT0HheojXcEePMzX7zOpM3I2U5bwYk
G41aF9U3nOKRasbJWuFxuZP6tDgRmAH+dEzq4+wi1KG1plXDvUkvKaxfGEXRv3CFB3n5bVh39R6g
yYM9qP8vvby0Oa/zfWrXaCF6aAwEG5A+aSlJo6gRnJZ9GY8fE9D2SZTEkAqfabvuqomNlbe3jPJm
NlE5T3nMF1ht9NOiDP9uCOLxg+c+diniRy8Lw7jqOCbPTZewgPcS2QoJPACpKK6QShiYtUvW601T
9vPVHlkmVzb7sSCX1b2VaoL7S+On6vp+i/R1ywLhNvrhAE8sGkW3bAQZWqngH9CL2ylMf/8nm7Wc
1u0KouK5JALcW2NS0Ft2WIEJPbhq1JVBtpDNr/oWDiyNGDcA0cTS8+kvTWtnl5znwBtfbiXUiLaY
tovhx9i6hkuHF+v9wK2XUUP6NE1Mun8G6c3SG3F4T4HpnrA1zP1xY4COUi0ffAMrhxPsIVrOw5jT
ws2L7P4Gv/kmISmKH49N3H6XQVcYsdXiHjXBBVeMPHuzPcykVOuny1g3Ba28DGgB0rgcWuxYaPgs
RkVhizlxOO+aGOM2r+lupdFQILoEEjNnnvDRzOwR1bRHqcyrgKVhWWSqvnYRKIrjy/+rZCh2kOeA
MzX/7s5KaMck1oq7sKYU2M03GuzJG2o1sTC1bGHhjFG37U+qFPX89bXMBKLua+ikWuBvQDV1HzaR
HuDyaHyqSeEWcstBFggHFVqy60VHUneIVO0kTk/d0kHxzt5eus1tezCt9ZyK5UjvcyUMDJuvjc9v
MDXKXFFCMsGhFD13dD0iGYUYsMKo8PyeR6a9H1QuW3q4FYx+DDiUBc/HenuT+EOVS15WtX2/mUfT
/J3erzO0p6AJGwuceQINsSdJEfRxKQbgR5qIQXmUgeJxxqCT4qDfoLoKNomXZQi8X4rBmTpbOgba
UYcnROG6pBP4TShqkcNh7X0ZlIFptpFcL4hsECniB60XBHv7zE9EwG0Qnt/4NbGdfxIDNqbtE9Qx
HS2tcWB6wpWENdWSdTegYx1v88Zon0/178uCRY+yihhqK7JfW3mNxwHyv1M6oPzONmMqbVPsyGCT
g116y6oJMJw2/Pk/U4UO1Upb6+s2sX9iHLzdncsXAMEByOj/3BnKimq2IEwd2wz3iH+Jfdl5C5Z4
1PG4LDjB2Ax1G9Z3hpyrAlDtkqrd+F3IZLM6H1dKqS0LP2LXqnjjxSYhdxEPMt2taWsUuKSlj/yu
s5TkFbebtnWFXp5b7pWq2ejLJDS6wNdLG2g3DJ9Y40xzv2qswHxo49VZrlHpI7mIRVBcH3NRmaDP
OnW18pVssVy3lhMcA8mcn0f01TDln0N9QqTlQ3DFGOzo1KWW0l9wgbIOo4C2D8qT10+cv7FtW1dv
rygNItElqfFlrZJ+kQckN+SW1CKRWo+3CGay3YndtgJLN8oNU9BCrqh4hIiu0kYffjYpLEYUEa2Q
nDvJWzdLIb2DZ2/85cg3Qs2CwlVoX0QPGC23f2I73VemgcZmvalwEQS3CalaF/x0InkzpKcKPbxc
mOMtO6jpttpGUYxrEXxy7E4ME2WvdJ5IwNTqhaeNtd/tM8YEXjazFolmBoChWYDk47zMRAa9ZTcP
F2ZCIji5sB7MXNOKha81Q8gyXHmviPS1IfDb04c5FBfCK1/glb0O/GFob1zatjSFNwG96SVQCbkq
r/TyOSGc9iLASIOfh4/54grgkQumAxrjxJhuY+x4nH04CQ3YLI0j8+kn0FjLiyCjtIsWCzg8ERT6
mXzIMIwTTciK+BovW552/cVJk7f/9eKD8z6spHme1tT2y3HW01CT0VbQ+W7mYekGQRzfHIhQ0HXJ
sM3OITQBNwoz9wxvsdGlkvjXG6VU0kLxtttinijh+Zc9AAC4dxqwnIWfcKkxKzfxiCNVpxqwyEIK
jwtU7FXRWje8XhSz0xmtKnoyxvv/iS/b0uqKc7VyzYwIBvEN05BYVx6FhNPqzP7m4QWEVAZPI/jE
buDMG9jRsoiOnGGnCiIrplryDYEqtySPELZKPvpR/rAIu3HedacHtp9c2RyL+/BlZkGVKhZxP+TF
b4bcsfPmLkeG7pZet+3bjhPFdeyZShcyYdZH5tKvKwflL9jgZAl8KKt8SE37DG+72KEkH8sNltku
HmFPZDuZA3nd81UrVo4fheJWR6JcC7aQzLB7a+rsQuBi5HLJGJeExjUOyStR1LBjVTyESykYxyew
9NddzLVTZF10RkGYFYRJlxf7dbHLolQa9YdaHxpdNGUqrkjyzeKYUbaD6t0XVAnrXS0DpYpWWaCe
tHayb44v3keKRx42UkpC0l6zlryv0edQX0YyBefobF5pm6C7SNZq7m5IhgH3Ewr14se3p0soWbqe
wjQhYqzTEs/0KGaAS4nQeBvO2kJ9v8LL8HokXFlMRJiU416WP2HPmiriLdztqPZLflYcApqwvbNg
CdBrRohco12VD6W02azdH35aBlO+YbEHhJQHJB2GZjmySgsouY6VmrmEz4bJF43bjdVS29vmcwVM
hYfaoE5BDsmOw9sK0jRODnAPBarkvwE4ra2KfQMJa5+k6NvX3+gOl/ZawmVtP3MrLmsmg04MuD+a
tzc10OY2DYxZsXENf7YKIJMRm+ZouurzOP0LgPM3Yw+F+sOpOhQla5b9wyz0+hqV9EuSIq0C9Hbn
Ytn9KEWTjPrvIt/z6o5gjh0cHs61UUyotWE1VBGwve9BK1alWcXzYvyvFIQDmhRoasmttim87nm7
EPeIPabL5g40FyQ+g5/9FoteJThRbD3RHmElQLC7xxr7Fzee8QskN9eL9AOw3RK5esS3EwPPBswc
wIZRIdXBh6eRvJB+Q6Vs55+DOgzJ4Dn0DNA1MwNxgmulGzLPAVWCMMGoJQ/1pVUZ4EfhiD/ybe+5
rkhgIqcWbmnC/tqNzoMeBdPnSiw89C9X+F7EyV1d4pJ2K+ma9DUGlqfPMfiYu/x3NyGsagBrFbzb
rJ7xPFw08u4oowiDnmFk3Z0cpdNdgrkAw9E9LOc/5UaGjRKoRpssc2nl8sz+9ffX1ix84CnIvA2C
leIlKJIclu4ZbwqG7aR5JpU8w6nRxR7b+Bc4+UTSojmlEPsgd3xIo5LLjkw+XSSXdOYP9qdQ7hrp
PmQZHCfT3r/mmcTzOHtkXah0IobN+wWdbr+EzO1cWzL0gd/f94kjuqENfvcVQiD9Q4nfIMAN5Mv9
/PqKTqKQBf6g/qkYS5JjSLR7ODAvBtGlwJzPUUvWNBX6nq+JxgZEhTRvHKpGOjxnWITXtBqAYq7b
pfEhBVlMDctpVOV9gtkbeNqTEt0A1DRdmP2bijHNAtYd5cBG5XbvUSOt+cttg/KmD4lXINeNKPUI
c/3Yaeqkp0LbCUVD/kHV2/NmIbwjCAzN9EzMQeqD1sjC85m6mi8lh9PVP79YWpvLnrEeyNxfU3lR
f7yV4nNsYeiVgPKdfgNgbgrtvETXD82IBS4JdocxP4/WApu3P8/f2R1EdhjFpUXaMPUTXScG8rlt
pgfiR8B1M3AkgeJ1Q6vwyxJGcDQWVTFRZTtlCYNXC+UW7A7E6CyspedlmNEljI6+BdaUZ4HDflQx
tSqXYzfv7fBZOttMJkP/Av+uJzXweyQ7El+5+7VBpZXBABNK1QmwaLwCjYiKMvoLU0+EHU7Z7kiA
8IVH3iLWd6SiQdA95R+cRckdH3gvwC37o5iQzBV7C8Wy7S2WUGsXAe5TNsIGI4RdCHQ73bOP+bCZ
Yl7V7gCKgNnaRFS/MxcW2Mys8c+jJB1ShJVc7NlSIvgu41EhLmXlzfd32RutebHKZz9/SYlYJaiC
Vxpa5608V1Hi+mrTDUKZd0zW4xqgQ3dZ/MJschzmx2W8k6Q2nkBXd5sdtXzfVdtN138AeB4h/A/1
lgY7pRRSyYadEH+9fOgk3kP8FtflQ3inHkgtviZroSeoRVBE5R9H+QoVq9pVR+pHuRYjmn14Mpv+
666BhSIoz/liwssrBpe3FiB2x0oYKE30DOpEsFj7MJmw1HQ+BB+PmQ/mMn3o06rYwiS0tCmQ4vLs
/zwpVTpgfqxXVwmVGK8RO3Hul2A2dn21ZXoYMjJntvxGQlOfElqiraWFjcUE0lot9wk5GZl+kL22
IfzFoOsONEgXqkLvSTs4K8UbiP/c6l4a5EquxFdARnasVUWoKBG6AabIyesiWZHodiuZyihNra13
h85FWCVBmPOwKqNbmZTxR2N2xw3ErJVMhoQuhe9+zotR97ubeTAiKE9vmueKTGarfaBogRM1zrDa
fYTDeI52NiHyK3qvdszHdASfJvN/YTB5Mwoo4INwmizjEKug97Npk2MvdyVDbg+6X8XBRQEDyYBg
1/ugtbw7lCojxjwGH4S2yOa42Q+hWaecm8MYdTSpvIs+1ysIR7+fa3NJQvOuPhX6x5Kr1hjxB/5V
XwdexoSqRxrMmM0LqKpcSohm3TVFIhaO0gI9YoqF63vU3RmWVAlpvKXU23bMhAbuTKPYuZm/UceM
LsLZBbWkblcUDoCWlBBb1CAXuTx4o/7QkL2HWu9c6LDIfFF+kkfDXuHZOFhiAr6WxUeN7Cg4IhwS
bODAt2I0YNcH+vTw9fW///5sMQ3SVCL1fjjZVBlAKh//6uEr/nOAe2KmET4kZfnpMdOYXLR/uIuW
lmHcFz/SnbTWIy87V6CztP8ZBhRJSgsdmypKPC/uDOEjZRbiEtGTcALqb6sMN8JuICYBOb0JHNbu
BKL3VJI4Z+iE8B46t3oX3sjFxzD1+RyQXaZgvGoNxbTgWDH1+DMARF91xCozf2vDw5eqpslFF69r
NwS6/io6+1kDe8fjMEYaX2qVG2PJzOPJ1OdrdioeZxd/+HRG62slHpVn2OCh+dOvTiKAixbloVOQ
EIQx45yX/AVE07KWHe1rGhy5yxB8/4uc5fbTz7n5x6z8SzJ2WZzTQrSd/6zm+Y5kP83pWmVX+Nao
ggln9shIVMSVAlAj8963IrtD63vgTlRi1oQDIq+O1QmzpvNBxpHbuOB2qVspqRSNAOQZiBkPVaRr
Uamj1eU/3J3jWIkFRom+/ExMWF/ll+RDsSIPfLa3kBDU2wEDL3RI6W+6q3r0EUnFBLTasKIm8G85
lTlKKbDZ8aM+H7qGZDXmk8oTJN6wVIwm7/je+ryR4e9tbIi5vCADPOGsOicOnDs9sg0dlm890Ew1
e4Gz2qSluxy1HOH7aay6VXscv19RAQ0xDxFePR0n1dY09O4UIL7XTdfd5gMLvoMTvSSN62sPlgHb
odvfJLecINSbQb3hWKkcMubG9xACupW6J3wbV1RL9dvHxqE3pzL0q/4XmpEp3+QKhKrdTZXxF/Kw
Q8Y8MGZdEf4AwDc5I6uo9J/OJIGgF+QzWG72RUaV2KTyXue7YVYbbO8/wpFTXTqD2Zkz19v0iHQE
GxnMX65wpJrdJ4zhUhsg/ftyre5sKfQqHamPmYJf4pWAM4qPDKHdxGBHJHgojAKqrfH5lJFFxWrc
MDYz87scDJOn2KrvNLEXKNj4nTTMrr7/2oI0SrtOzwCfr9qdzNTB+wS3I1/+hl69WpC3n1tcekFU
df3CDbxlCb+AvDNvt5rCstY6P2V5QzmsaX86cZLI0uJypcD6mNg0ds06b9RAkVezH0GwKOUcV71t
ke0+ndMgE57dJdCUluPYS1zlrFcpw/qJIVYa62tHv6IMUZN7cAKjzUOmoLUcI9rRXKeFz9cHU3Qx
VsGMnuA6PE0524ShgGw3BKexqv+pNUxaprkMtylIHjGp0BY6ZEWvCSvg3s0ek8N+1wBMLFiAQ1lz
UEF3tIYLOFrcCGXqc99DMh74SdIB4pXF8RG3OVqD/8tVlrlOeFTxw1R6ftzvWu5BmSC7Riy+sXYc
mj9fkRj6EYdXv61nup6m9CCAElnsz5KBun4jdCY+a7dCny++/SwFaMWO+6dwQVi9ilH6I1yu0RTP
L2jNvm+XbiepWxLLGK5VDeMlIZ5j+kGR9VNuDPB9yO2dASh1gMa+c8E0ofrSy2KVTN1Q9EuYR50K
O10hkjlHT2mWF5w0TLKpRWR47RlrRl0QhISn8WbbVe6ORgNfoSjl5EmxguZex47tc/HL5hv4EyiO
/fYMg9qpePJb/Zril16DIZ0jWfjZhzUZRg3w8ySdWga22EhOpkMQrVibas+dDLWN/5N2nv63AHkj
xdxPeLcVcAG7VSNjfUW9PBPdfI5r7i9v49AKdGIrzBS42fSahDzacv7nUzM8iCvO91fFhTzoQm72
a21awU3OQfMxF+/0xtIXs9ELCHtbj8EzLRoEggfmJEGlQ66WRLBrIu/fI/TddcMxqGCOqrl6SpA/
kckVj8mIXyFWZasezakgSCm0kD5R5uqMOVyrTah0gWUxQTaEkdlCxEUkIgbhWLQD1J7R/Tsjaq+K
quwXzlk+xOlB5ppFPY5jrqcDd+JBIxXkT7UfYt0Gue1SxvjgHB6hgjW9aM1FqAmWAIL3yyLMuvX9
7B2XvL8Sx30A9kM6LDQvvQYSEYyNM/HCLeVwyluqUIR5h59wbzjmyvTnUkXDz5Zl4WWW7W1TdecE
3x1mSMkmgx3BdYelekOk5fwk9MYjLkLAwwpFnAhgYhsjF++ZQxjj8LCMskpm+jyxtdkCMhgDgdfs
GXXNKRRmiuYnRGTVUmZX3e8ojzKsAg9KopI9Kav4IP4fwMkSZQG1dKycLVleSTC+Y92BULTccDGC
LCbwrbAMuRnNAMtc4sbFcl1VGqe7X+MuSK9cqZm99irjp4FrqFilQokXDs+RZKXKb6pS94GIb2HO
KWV1xHtrpyniz3oDakxXj1mXF/GRM0O2J6iLxMuw78f2S0cN/VbgV25tJn5BekpOHf/qjtWvZICp
eAn9/AhgQNXPU08xtU/brL7AVcavuospV8d0LaTFcRxeQtSMPkLBKMmb5ecXoljQVuyNflkIuSTw
mKynap1byKXRU5sm/EIvp0sQivc875NaOFCZZalpiwb9FsIYPX8z+TDUmsrXJGM5+E2+3kOAxPym
7jEdYq6UO7LEnLrynJcjUDwqJq1d8pSXA6iI1Md528pe2rztrHmsG6q6AroYMO4JCuIKbP9pnacP
tNNzomu3H6QzhzajEMZnT4bk2Q0BObEVmPUFTH59pB+vMQqBRta/V49edtCEONxLyjxiEijc8SCg
Y1CswyTubvFNmjSocfStVStMzyXqRHOfyJqGH1pHaMx1YMP3uGsGuDN/WIo3APJYaqX4vSIz+hFh
fKZKT/rVRGoRmowN5gUu2t2pqSQFZmlXVBqcSHmWH3Tg/UTfdBm0+dI77o8syLfShaDxbeAtkmTB
THRWL8ot5UgOVkB1Tsva82VslKjJ/n9JsRBQkB9hA+f7MrpPNfN45N+trgxyd22HGtKcigSdmgYj
6AY70/lHXd4IdCWVEmQRE8ZqD1vGbBvmC+K2Kkfl5IlbCgRF0+Qw4HRRnv/SanqWgD6Se/frY9n0
2vY46oYV6P2PBYkyKaQjXKjzpXi4eMk9+Az0rxntaw6GKBObGaYnatg9WcCvj3v/HKbYQq+8Xtx7
9HEVxAD4wkZ93GTvhMlo12gvUKg4irkmW9SGSs9Fa+ASurK1LLaAlAvJ9KrVW06+4JVAycQat337
67cTrBYpNUmdtTiDkn4xQuS2mYlXDDnmd3OhpuaESJ7qKWbqCx3GUkEIHR9MFs/rGtJ+H1XgI8YE
vTj+x/j6cYy6OCrh+XFR0NG3wWPDggaHmvNjnrNSBnqh2KlAfS/w6cNrJFny39IaDtUMU2CbJlAI
lodFuhF5KOqV3iwJWtopFyiix7mX1bRyH+0S/67AUeYImTvmy8CYiuEzd/BnOZ7OAI3PKMUfIWuR
0NfP8h+1ImOkExs7cO8ZanXR0mLzVmg0T1yM9zfxLSvpUgikA3dccuvTQ4QH5kZx3NbQmr3A3IOp
iLLYmgefZoSkF7x1uWf9GEE+Ox0ffNRwSQ1X0DLQntndll94241kIoxDQkPeVXmUH63sRhXcSrNh
jdcp5SKXzxKUSmE0vPGgGsMcrDLkGmQNuEl5weULIPSMbJtnEbdaGHLuI6/5Yb2FQw6k2wOMd6Bv
MJu3NLMSUqW4b3AJu1kHF8lhU88uk5pdbVok9/mLZnLTPAiHQJXdqzcmECAyf9rpnjcYnF8c0+mV
M4MxwtZpaCYHdmz1sXsUhOMOvMzx51E5HCB53kTb4gPh1hOslGS0qNmsAO7fd1bJZAsOs03so6u6
x/pQzCa+dS2mbu2eJQHfEbTNex9XnBAKjU7sJiuyBLAzV+zUx54Ff3Gk1c+XAvvW1RqiYa2uTpTs
+H7Oi/6ZsrjOXBNsGIXQ7GCIEpSV8AdPc/vlYVdpH0UKf9O7guHnmHmR+4DBHojSGbTIYB54gw7A
yu2RUtiYGizcijZXOChrTkfX0tgWDJYkqpDa1/asEK4GYl3N7A7Jev9BEfSgIqWhHTMiAhQZ4CvO
6lMhbZTlwkSgYjvcc3Q4A53ORHsgyMPIcc6+XUcbpXzh2kMw1O8af+yRn36rZxSnQq2M5AtLfwux
VEGBDpie96lQTfS9REOJschSKmB6jxu8fOFSTFywMGlMya6ucVWuXQmiAKnHulpNyowTMy957GI8
cm5Y2HS0MX2EJKUfjm8LnPIuHbmF+8VLWQU8XW7wIjrjcUbJ3ih5GFYLywjrD28kciCPCeCUMTSU
Pr3Wy/Vcwob/5HR+2tKL68LHEjVx99jt8ITlatUShXbEjse8otBjy9Z5i9/OB4XZol3l5tDal213
/pv5aMlwrdL5cSy1avALiR/BXy2NoO3jUpukiBCXw/lNE5SUXrFS8j2de1KgAPzm/A2SZS8lN1H8
FAkLNMTzHlo4VQpGcunku3sVt7njsdnLxHK//9hvq27WIbCJwwBk0Nwl5cxPi7WmbNJyR222om6H
xrhdyoMYl6zJ+p/Dd5N+cZa0Fk56SlGVWHNFlu9aFzf7lqB7ReIWAssXnNUCIPXYtBUGssjULXHM
dHQIIs0cUpmtcJRX+Gwwus17IlxxX5L7tLPL3+Dk84mM8y5aLsmPqFvVf83ZdIsO5GMoRljk1CDG
GNZZaKTz5IJ2V+LBVZmiV3XsECAXDa0C0lVzw4SspeDh7lW4XyCKgOZZB1+S8LwS3bzPAoshMzEY
I9R8hAm/Axa+DJKtHqIRSufNOXjv9Lv2F3JviCYbIiK3tz63AQVkjkoEQ/TOJiEsYBPUDGo9CFuB
PRpEvUuvO5pZOADwxn7RI08/17H1XIJpuW2Pt7rIzMl1WOB2qaQ+Ly1jzRXU/jvpjgFIzjw9uOZx
mOX4wLoV+/QntUjtndTMIsKtzzhC8B8CbOY5OOBSkTjVBmAP8ZmxFaTKhbodLwkGUYINXJYemjnN
n+JM0UagzERmo9lvenpFsX49C0ulxZoIH5WUwQrD4bLOcm/DqjWNyBfIlsTZPjrHkdIqWV+xtI6m
QoRfA4d3az5pHUuiqorpgIjH1G0gcJalwhJXeLQK/kujVdTieIUG7LDppnFrwbEYN4x5J92/xx6A
QnmIwrb+UI6jxH1BwMeO6VemuHdpz1pHvTSeP7SEtRxW6+uamr4KC3StTNyq8xiFr+Z6dsU02z7H
WIn08EHskigvFDu9KWNrON/Z93ZxL2rubm13qlyF+litr5uYRgt0hsowEIOObwJ8G5gFV3OHnpUO
UXfZtamL3ioen8gI2Dn01Kosw5V24SAWnXqMKvRSsM46DHQI9OHVmNXbOsUt67EI6BNS2rDvrYpy
bxySxDZsxjETi1jUP+JYspwfZg9ya+VQ5iKY+fH1NpERSc4keMVoKruO0uMyXk0dLkRnE5dogEEf
cm6LIu2xrfLDjEVyQSW5+Y8Q0rHiJ+MdzqgU7jZqKSaLnz0u3jILAJRsGXSaQreJobH8d8GoJcSG
AeFBBY7lRyjSgc/6JtlaqK1xzHeZnZecVswooy+lMAJ5/czNCOgSOvn+Ljmvb9aPSNNfWztX/dLr
uKr5Il/uAuLROtxKh15KamF4z//sdDwCLawzTehbigWzv+MOoVUzQIXtcm77MpDxMFcsRa9F8Tk6
B4YiHEHQDC2wjiNtxhI5N2iN+WfP7Kunf5Ni1oSBL/oWfiVpBFFcn1ZgLiu9xYzjt9LZvpQ8aJkl
rbPpvW7WAtI8d9Khwx2lyvAcdySFiCXvgZBKgsR6fdXvtr4xqwl5JNefF7HPbhzfg3X1rppx6QD1
KzYy4dxUCXg3yA3LQoMM9kGjs5tzvnC+fAoxt2bs4f5Z9T4e8/HqsjzJgA8S90vZl3avNStlyiDK
oWMASVviYRdupnZoDbaZizolOtb4qZ4I10uf9Pf+BUNA4MV1Yuw0dbWb7wSNjkktsOkc5ZfLmJXF
WMRP9J3s1hSc4vUqWWifIsB5HGALXnoLhCcrKuOb7wdXsUWrfyYnoV7tN0tJuYxAt5t3X+t7v/+5
lm90xuo0FtJqUIkEEVQdgGwX3YCqWdi3xDVxShyYog1wTEBIBQeFJURBrJFlBkEaU2Ms/GNuYgsT
ip4e/sRVFAfi0521KkwM5JdlO6JmOmT2imk+40LJg4PPvZRwcsNAtMj5EX9iraGA+7vw2TTaUaHd
h1uEAQhoJFh4pcs+qQE6JZ1wTC1l+RiTNKOUtDKfMPSFugU+vDK10wXf+LQrXuPP42KMxtuu/Tnk
eOgTvDig0EmzTaC9UO98DQtEHXUY1arN4zOLE8XQTfmwvOs4U4X8ppRfd157x/jEk83zfYlvIh72
W8uezXmBbe8uHb3may5+DnQuXcq4nA43f0B0UVtYYv4ntp2wnyjV5ZHeQYG47pePzsh+fOtaSsIj
V6bJ9kfFbv5Zx8i4LMH8Ig8aFJH3Aqhp9I5dnR8rzXgVdKg9ZxmtoxYcunbhSqjz2oVGMaYnkN7d
VGil7fpp6PhJ4CuTifUr2ByL6/xVCeBZdoMy8w+f5vt3RYBoy4MrEkq34wh7X0F/lBOIstqJ2vFg
lQUCMiB6gAWHK3wVCWcPwlseZCvaTFKPMUdQDPBSgWNN3+aQIh0sjd4ngTU82eHiZAWa5Ybv81H8
dxES43eavhWdO7LhLeN7RigRLKKgZWqgQwgr4tpjvOkD6oEiGxjoL5gnGqH/93BBukzHneli5RFf
KbdN849NpHePE0E/QnUS9ZgPs6L3tkTtjPcCZbJvDcUpkE0rMp2jVRa7nVSLfrX4L5VvUKHa7npk
WQpyxMNpcQJgUSyR+ovmz5HDow/Lo1gLbRTiWi8bzOzIOB4yrG3+QJ50uzb6KElAqkeX1jRijq0y
0/nPTXq7ioBdnom7zFBgEzVd4MsqUGZSnwpkqhRR0cqMBZyo1TK+ZGwArS3/PXZxVtfa8d8/jypQ
WWPJK9gjCMnThRonImylo/1AFf2xGCIYYu/CdNkOUp79KtVeqQv9/73Ge5lnlvyj1GjJgdpFi5Kb
Ymo8uVXcwNM+IhTGTjD+0dJg1B6ObhVotVgq89y1XcuiP4qrAzbkXYBgA9dLMXS2j6FZPPSRhinn
azI6MP0epZxQH5V1tY9QHuk0gb+BO/T2oDD+PIX7D7pmKPaMdayGsqbi/V7AiSJvVlXrGcZmjYU2
wKU3dH4KjC3iaQWpjkfyicII3hfn8dgIGkoozC6Qo0N5opK8863HqOm4cAVnUDLlZR3ME3LT7wKc
ulHACl2wmC+usT7nDQsaBLmWFggcBerugIml+PrB8HmxhyDxsyfycb/cR0CsLYZbM8BrGo1tVR8O
Sw9orGFk0cAc6+KP09e7svoCL8MJvho5hu+Er5zkEH1hJp6NiP2lNYoSVtLGD20NykZXC8YUp2bj
orjKIRoA5r3Z5iHnv8sLlblTn0SzAFEcrprFH/X+JR+/Ih8ZpwNxYCBkWBxhZAoEhZilH1sC6UG+
C/TbEBC479pXSaRZMt2ZWUiHYxOuA6QZa1qIoy3TVa4865b8GI5aFLloBnkJHJSGk/Z1U7tpxt+Z
iWRvHvZu3b7s5vcB8Y8v9t9JNNmznRpvlNAJJAU12bVBzOwbmXQQSBe17effVZJRM0JQpVw7CVTn
iocb6z+R8ThPZS7gcL1vB+RDahww5h1Iocch9gqzqH1B2GEbMmzmpLlYr6J10D0WF/YcAZ6MpcAP
KkEW20IoikjSsvW600b+E6ZepstDYDNLl7GiZu8PZkNaNOFE5QQGU55eHG0jl/DzB0dX9hxib6RQ
N/QTujEOz3l/Tj90+mURi4ypMSga+aMoF6RnveF/7mvSPTy81E7C4J49voaXXuemGgFbhnXrNhk4
zfMb7/4oTje1t5c3y6z7/QTF1nHDJw4NCRg0XcAcLmUZOeLYwIYavMHdYZmdL3QmA0XchyOQQKjk
wTDN9IxFPbTLiKcKeHWCcHAUT2wcWNIJq/4Rly68cfQLf4BxqCHYZU1aF38aYnV6jjeIvilxI11g
wN+YJnLBMUHRD461jx3jUOddTdN8wjllMfjQOaJz9wVMHQDOP1R0CZqarLL85HS/hk13VLuvkcNq
Pw8UCJzxli6jiDcWfppBBYJkTDFcU48QYEyzpBnMunVQZqOGT74VDNlga/+8OsLi01QaYDQCkBgu
248qaUGhavpSux9kz6FtavbnXEypnrGFnS/Tnj6BBF+3KF88MSQ33jjqztp275KwG0MtYjv8f2bI
YWzd8qJtughyDSQhhA6cg7OMjHN3zRL4/lV0X35URuS8QppZZJmeNOHg9AO1/vu7KeWWg5DafTfY
JXH0BvO+VOIi7nWjKdkpE4LNyL5Kll3jC62KLjvwu6VRJejry7VNr2x39u0P4XxsI3MxRfzp1S3L
1gG/a8WXDck7/KI5lbYg9dn9ZjDn7wYd9wWbMn0TpSxG+yzebuxm2ZyOzf+GI/nWKyzDm4va5H3U
cPKHhhv+otYxDgWalhG5YAzxKCHmoM4CLnHoCEGdhMEXWDY4Z5U150D0mdq55XDCQX0kgcu58xPi
yLQZzjbpNfiaa8ycUC6QUclqfcb0v+wf4Wu9D3wY8/iktDJxht+lnMT+fIVsiLdbIhZNu83uci8d
RmRDsvfQ/RI8Sk7PbLnaMCkzTS57LtIsRUitjQDpFZwWvzXNj/nPbcQ4QrdWTdHwhr+0jwxNcUYA
y8RJ+3UOhgGgEGwRboRpJfU2SL6M7LSN+My7f36VHi1fmvHtibSzWX44DIB1vXjufEZx95Bse3Bi
9pfgrk6uMu1stiq9EM0f/5eBa+cFdqYDlo3YU07/Mio6xo/gTo3hiMiN4UR28t3OMdV7DeQDZewk
DMxtPWR5KN/pO9qRYhd8o7Il8t+6vNTsZexxvIZR3wVNQEEuE+r44lV9te3AUA3rDOiFMoj0rO2/
dm4jLuH9kipFyvmd6Id9Yr0LgVJSAnlNVNnDgg88POpEKAZYdC9/OPgzqohHa9LBr1KHwe4POUVE
mjL8DJWnfrpZgRBNxykAVl/l6Q55z0FE2FY7Ann+n26KI0oYKxcIRwsg0Xd6uBG/z1mVNlXjQVlp
K/zaJxN7BcCMrN0XBR1Lu7iqJDuLcl3SH9WrZ++Ng4LvNwnwzeH0hfdVuDym9zpfiShUrNJ1cxWA
9YDAozGFyuAJgDrnma8p8y1m1tji6QDLu4qKkGMjCDxNbTN62VnUzPdlGNYutN6xY6pmGXTby2eX
U5aj2qeyQruvpylFimi9odzprICLwsiIQrpYtkI43ug9P4yKbzhqKcv2IUC+MDgG2vGiCvYroeBe
WQQ3JhT+OiaaorgNrnEDSP1C3b5AOw34TxIqJo3s+OCrUg/3u2yvfGyAjik0r0/ng1UM+aVUS6CC
wwCdAoVUOYq4cxAQfFsM8O9fKRMMl5m4Y2N9d5A4CBj8wMRR1bhLauZ5deFnI46UtovW7se9DdbN
S1ymSjU00yVEXYrp+i2avDx5gnrBRxGkLsPkRsjkRX8KtkidEyW1sa+FlCDnc9W/v6zlkE8e45o8
GRzhDMlbejbfIPJd7ooB2svX6YSFKPjI63qUxda2qsWvooS+qubs5nUfjQcoAMoBvXrIbC+K+4y4
wcVZGY9U4+0kAxbA/4UD/zS+dLj2heazuR33MO4F8yW0BconmPJe6Y3stz2jaFR4CRefcHbr0nDk
x/nNf3+42ijl3DjxlUb/Ei5NlWaHgr6l1ckAR0y+vtGnmGWmbPnE2Z/ooa2niN0W1nEH/+Rx2ycu
GXDRPnZatKT6Qwe+t/1LulFGp/pElGreHjbFckwc6CndaCPQjFquiLIutBqngLxQ+dU8ikeU0xfH
7v8V2oh/FgCxYuhzRrs3QiuMuChmZgtvMRVG6Vp/pBU8Jewik3DsLN2avLU1c1TlocdreGOBinht
pWXFDhRqRxyJ3J8GH8AckIRDhaZDaPxTtRztTf75CPNVjKnVQR4e9SWPCTE/tsWA2nfZghyN1YXR
rOMZf4ZXHhiPOpm9LfrK7cQV5kQBOwclTWPSuUuoUEhH628Y1PGL4fI6Nk4F5VxsM+QgguySBtfS
MyIbcXPQrGBHZbY771ZDSy/opdCSOWumi3TVg3BzaIiYPZnu33pgoQsAzTj+7FWYeaFT+Liglu1u
B7liVea9wEgSsp6NUiQYciHIMvVjpgCdgfRPVFfNts8QIKrE+aGJAwYS8HgI/BGXCzi5lIkVtD5q
vKkRQpl3ARGPAdnpfO6b6ghFUYou9LwkB58Nfze1AdU5UgSyL98V4RwPkj7I5Ktd+53om9+KhizU
ILJm/0s1VG8Ol6jJg93TKn3wEsotsfBnAa33yE3nXYmnEHGtuOUpjqkdlJueTk5Bys+0HwL3Hwl4
aJV5zbynPzw8+8hgyzu8YjCFeYJMSNTjXW8u3xqmAF6o4HXhAlfgzUEPQQyq8RzON4L1rO4iGcC/
RgRnAHRuubK/D6atFJf4lr1gxNol34b8Kskytu0fY9fYY5yFQPc9edCKm6QH/hmhO5810RONAn8q
lKmTKOtb5tBC2R/i5/5qbdMpiOqc/mdWONKSX6k2K4fiqDeb9aTk4RqEGrfCjvnrt5kb5uxLKGt+
PMazsvD5PJUI9U3lnq7KyBGshonWSitT+olg0rMyAzs07fgWMloGY3wKDOuRG/KKxg2tq5WVx7sT
MbOOJYfgqkoYGLw/jucuSbcX8LvrZBYHrg6gCNBmCkQVGrn0w1J5UyedmgW5OOup8yuOj9bS2b/w
cdsHmbxF44V2+KJJ/P+UjffyHlI8KN3vIkuc/5OwjDpNc/jg6QJbxK/LE3ybwCmi9JKhxFwBTNlg
dYdwxlTjWBAT7I1iCHUkOrsbNyR6eNcR2Wyf9S7fvnqdnt6QWSg0TRREjxhQGuLdAlaHNE20X9/E
bfIeiEgJ+swrInKLzwifvDXaN0FiYewONTVoMAngpo3oroUZdinu1xrf21RtAzJmmr8DXMdvRbQj
xUa1B6+Eft9cLVMfpIgazGbZz57rb8rimJEVcymsViFIOBsoubM66IG+DQQO+b64GpULBGQuopW9
Rh4uenYWGmwupXL8FZ5q/v7R2H++fevRlQjDO2nXVbaszMo1DqIfBfTG6pp2ouy3NG+gZx0kervv
fHNthr/9lHZ4WQ488hZO2bDbxfF9Ef5WxybQpaK3RVT0LNu0Xv1PwRvS8E1FttEYDykYPmqmbWfn
AN5KD21Glp5YRRdZCxCBdQsq11IifhP7MotHposw6O1WS0vCbcAGHsCDj3w2cWw5qiLIJXaOC5oO
kNTRkPeWrk8DWzmYtiOWD05ViIowY/QlphqB/AssdoBiXzeeugdHvTCbGOGd78M9d1keSszpVKwp
IZX8J7cOFVHhsMQeC+MTCLneX5vrV36uGTsPl49PcA/7m6JKkaVWpk3qjbKmLytON/d9jz9pKkTf
Oh79TubhVrNdNmH5YPvQBA3+m1eXSDwdF9/ejt8FoBDi5TP+uIltZb++PUBR0XkCLyd2aatjsHp2
0fEbo14IwJducWlfizmlJNeqPJWCF/B17eIwGSf4TLHUCfMk4EUf1Bu3oYafmIFtyE/KkUyANV8v
XCLhrKtAqrkCOJ3V8tAVKO1Z55bZRgiUBSKe73ZcQJa5tsZ0Wtp+XCveNvyzo86GALIFUHbK9pnn
LwtCq+xheoAo32J/rRfEgLzVnXlmZWHZt0CJZtNL3bCpW6OlD8o4HWFcBmRVAIcST8eKnsr84gPZ
DWgqbsj9iO6TzZkoTeQ6eX2Ga9/xlSQGbXSmrvkGSp4markIe50NIgbqQ+5nd5+NKhajOuC1WTvx
9Bkci8HE8YDfGGLhZHjmlZbmmt9UoeAZXmnTkOydPD+fXPdTv9TN8Jqyh/KQNgxyxgPN4LmMYJGG
IAR69+kokQxD4eZiFeSnYzSmRuUgDrk5JiNeTkxkke5DkwdRZveJeM2RNDRTISrY7BaqCzqfXbl7
zNg//8+rStareeOq1/v/EFodxYlseDOBt9ulKNI0S92R1VjlY3qe9GLewlcsCOVkPiXfb2jRQ6tT
l4ESqyiVlLzSL4rujPUhnei+LV9BTZuwmyyCORdFxw9kV57b9x6Aq77DcYcId6hKVNOJXpzUH2F4
ysN5iHXojnbdGv0qEP/qofcbaiPmM+moZUCmRgIpSjtQRdI360apm+TLipUgmvDbkawivnUrgFf6
rR95hXgx839KMdyOS8IQ42URGWGkQnGeYFURSXqEt0Joyj9yELdT+f03FFo3xENSJjW7zn3c15tf
r/7DhnT0NmNhONCay7BkdyEcVhHjnVkPoOFmudNWnEmXZPIVAbeZ6Gh+i0froOaRhO7i1/GrS7PJ
F9T0VpvFVmrLP3rM3tAaROK3Kt0vxbxpSc6ceWfQeFQJZldl0dD7MLewe1voFxRD2h5307sTBTOp
dSGZ6bzx8clbRSw0PFYddXaeH/oxTPoKzqdzu/Nq4PbegJ0yHRWILrUwxgtO7uUUH8zyeS9F0tNa
po9PuiTHDfYHMG/XUlBoSsUum9d/TawetiY8kn2lbVedQ2lq/4CiKqP8wWyuxqBuN6hZ7s/dKwte
nAPiKQ/XoazlxITKbfbD9qMvBBIAfFKFkVJnCYMpJOnI2SipjU5SD/PkZlvxA6LO72tQr3vNN8IT
c12TIM6ujK2NWdrJPTF+qUv8QVKpksooNJouNgMmyUjMvULho/3chcX5bIxftpSSIFBGKIFCn6HX
hJPMkQsOhlyEKrClEaIFS4dmgsOt/YDH7e0RvtdSmRT5IqSZV20ADLsljzPrPJAcwIK40D3X5+80
3rOVB8cg9VpnEl+dJDnGaqPVIuXatRXoEifdwFNbbNmbuyiRAVNV51T8Pi1MSZIIRqlHQdt9Vzzp
yHrf6uEZ0lMZB+ob+uFz+4yx7ACaOtVd4vBHvL6U4R/29PlRMbWQvb32S7RsI7gOTxbxRREpZEMc
Cb82+tEQpmOkdV6rruvi6oAJB9CbCMth27aauhte0jeyZD7G3BfxFxl6DJws0mDXge1fIegnRA+B
qLJTephbg9oc6VDowXsNBfHajjS44a4FxJOL0CwJ3aj4Z3+pcw/HVpvIOlfqpoC0noEMiflgLgyN
Yho+zrAsIwFgKQ2ZYIh+yV2ElgWfZKq+06jUSNbMtozUGIT1zlAbv8R6glctvPWLgeyxliW7wFnB
ij2/AopyV7oLJ1muQ2fDL2SyVbqwTQajYImhj4Zi7qUkTmMdscPPnHJcSV31PzfGTKEaA2j7H4/A
8XJWVWl4wEBeyc4GV6JtAMxlcp1Clml+ZHRiaUXbgKa/Ho0ZzS1uvAenfXaGNkPm0GdKgq8GKQbO
BJR/sgtdc+P4OoXOgeGuruAREBx/Ak/Ab023cw/v6Nk5EsqeJwY56rx4Y1s9RCuZxZeDzidHXs2J
EkPvz2aotY54uNp4vVvaAiEeHP08+tM1j80tUc12hsaWKvYY9LMf0MC0QAXKM2F+lR3PIaS2gWoB
Dfi4eXA4IbYnTDXKpmUr7XAMxNiPSHr2NKdYugPL73s2xRPh4jzNy/ga3yyhDAJjqj30vlpHGl+l
s6BIJ6WTQfyaj3IS2z3ZEYNSpmzhYDUbUw1n0yZd9QoDdy+ICOpT/aRRH43DpS4OjV6D+qHVc8Dd
6DeWBv5qSErX3DgTQwJQo6XIigvRavao3T3sT00nnVBAbl4NhZU+42mqJ9DGYA7GRQfHC+JHu80I
4EmbG+HdBu/YmsYrAzYKbRZTBNWAJ7bjQsDVnq80OkNhBgEHy1HJtW914z8nFQesiXgl2xQZ/OM7
ixn2iQ2vOoq694S6o0TXDKamN3yTwi9gDeWa063bTt9IImHhKa5OCJTq7ASwvB0+BG4izjPFeTkR
5sBVBBk3ClY7qPrlS5PXv3BVFdb9AoHWndVGNMhooDKMm45HTo5L3skJrXWXjbEAdXZw/x3t+KQd
hDHBN404CzqeXc5KPdCKx6g6TTaOWvEwg3WLUnIURNA8+C2neWh2EhZPIL5pbFd0l3gSuvAxKOUZ
AAtC4csiOSCiLN3Jey1H2DSHRkFNSI8nKeOV7rqJgTMFBeKSSepCthk1ZypqNG8nmz9f9rXzizld
Efb82cV840OgSjQzggMrU2hKNLbZkhWRDK4ovFrgcfhQa9IXNyhfKQnozKZth6FsFSo6nu27PhxE
FEZvabEuj9MvwcZIOHKGPXGtI7jQy+XvpRhu3oW3LZJ0wPvVsnWCr98a7daf2RMe/54OHcn/+d5e
Zv6Suzfq+FSPa7VjDwHo9oUah7VCL+TxjiKmoa9xlZbtrFqOLpuCScPOQKKkm7QuNE7sq3Oag5yk
5gypJTDw/hgwrQkeehaN/Pl7ML59L33bYVvBHHpSBVRSAOgyzpLUxmuAq5muyhqzSkPIj7vXqhw3
dlxisj095CH4FzLtoWg9aQA2XmDoyV0rDbW0GqDtpDirHXplcQ2HFgUyNU22GD35PNYKVWIEHGCG
PoFwIYZk6Go+Yg+rU8GKUPgbUi9AWz4cD8i2DMCSkKvKcrmWyWTMbPuXukQGjjtdjvSoXWzxE2Q0
diEFx8Rtu96ZHNq7Xt0qBEzo0JGC0FLyIxsSNQ20iEJM92KMkwUEjGTB5FdQxglXzt4+c62cx6HF
EyOiwIBW+PPGs1pqzeMU+trGrXPErw9ZNsKXViuluQqwQC+EOlgTeSyjSitGwG1RsRsbzLNFnIz3
RYsch1sz6q2QiOyUUZhqzYB7wxoAGjowB+Xk9K5oK4iE9g3r79tBpRLipdJI8Cyd8CUE3NKRaEES
Pf8HWLJ8UelPrX+hZ2OPwmugqdpEIMNBb0XbRWGjTLcun5myPWKBymRvW8stDve/BL+ndwLsK6te
yIvZOUaiLwYmj7GbYO7N9BmpLCQusrIYiTErdQURBViArCuUI1vP/G6giOAotNi5pyCM/dIrVoKw
v1Z23Gz3ACPHaFzSVkC3GpG1k7cwG4oCLVTBI8jk96rNAoU3Dmoo9NE7YgTt8w4XaiLJUqNc2gHd
T+JT/XL2vRL7q/O6KiiByyQUJ34iN10onqG/UCoVPU6pzohpqjaXNH5X4UgP7NOVDukYFVdv3hiY
CRvzqhtrcWiffttmCWhJR9YRH1u3TliVW3byZ1HiXbvKdH8/lhmIfUNfSNXTc8LIwMkNMcMpyUt3
KEbGip3J6kR/uKHi+qjeNXGxkwZgdap6vpjzgm1zrtwELjRRSmepjafndbFnccTNsn7Mhatl/a7B
6sKpR/s9I5u+UId7hgQu58BqCC0FXLTGiEoJpTSG1dgzQah9sOe+yEIJ+4/1ocSwY4j5xUl95p8p
tDN//rQrTG0uIIgmMKabUeavWWkup7sCWMaXa3KRPuxgT+3WEC28J0jJkR3qYn9ABb5qvUXIBuMI
T10k4mEzaqxG2aSXORqFKoXrRhexA1XbtYHYAaQUd4qlY8pMeBHKTSo2873pyAbIH2QDR8QYK/JN
LPIeo8JcxIiKmSAoCANBC9UwC4YWX2dKd9z++kU2CLxJu0fBwT1pnWAC9hv/0SbjDiekCj7KTgjy
ypxrN46OqNq7fwS3N0+WADyBWQM/txvHarR35ZqcVfZp72wWGhEMkPteieLItKr0JU3aTQVVBgAc
srnpuP8E8I9tLmnXLO2xJwqCY6Q+1N+oJPz8OKZHa3hgUG2jhc2sNvOvwqS+uiW4KD8PWRAYsrfI
SigRfYd8ugao0wVuGPkyu40EjZpyJL1U/7sJwrZqGbuvqZVn/C2+DS6FM2jeaSgN6AVqHkvpVSPM
8C6+uYM+jl+TBkvQItSQg2tkCQOjshY2LRG5JO4Wqq7/f7CCdXtzZPI+6oJZLMM5A5wgdWnl+0vk
BdLxkw2LXy2V/4SnKC3ksPw4PNzY8SrlabHjJijD8ttbWSTiSzdJgWlhEXr58xm+USi2n68fo0TQ
Cp8Ryw/kNw4IvtrC1UYZXcUL0QcqWAx1jS8zSuoyPVyumWp0ByLXXf0CJGEqthtej5l3px3II066
ZasAksdSffQB8dSo7Iql5cUKFaZmP7SesnZb4mNNi073kkseVtSoYQRj4/c4qq0aANqWk2LnDTlD
R9A53udEmH2f0YzDziodrrZjGx2D1QOCNw2tc277dEcMdYrHFBN6QXv76f9eFcxLVNwPvF1FGOrk
C51g2/y9SvUTm9+3JgEoktV/xDSqeilgCS8ezyUNq656f4GRlzJFM5w3hvDPyU//G8Sx2flzzmfw
VixwycGIDmNV5sqNxtJwKfp459C0kU5287/KneZ1OJ6GZ9W/CgD2a5c5O8FEoULDniR4ptvKhZEA
DsnfBD46K1QbnJfhfLt4Gvuiiu+h81UdPSDb4rJz54eM2mcKsXHJE/5TWshO8OFgvJkJoCvBBx1n
2oeXFB3Kou/9QuY++GXHYx88S1wk4sHktTRrsQdf8P28yLL23XQhQY4aDv3Q038V6Fxldafy+Bvy
iu1C0y1VYPPUBkljDU5FXG+Onn2T8KEHf6GFozHyAkgjJek5Hy77UEIGhNEQcUTO7U6gwVbNS8sj
QrPLcNb0J0DbOTKFMTNhCQi8W9HBH3EmEdyfBJKvJ+RZPL1gjtwg3QXdpcqdd3fVd7mT5+nRnhBu
HWPmefE07V0GPtlRK5ocNxtADmByrVfSdTpzIv+XdBf4EzJOU2tM3GP9WjuzmG52CYMclL66UfZ3
qLCqH/91tZVJUk3SSARb+VYoKmZjqfPg2nTy1ZISITs9ZUFv2vjLP0U00V/iGFBnafMeFENviXrJ
C/eB6+g4n2kQIm+MkbsATioIx5rbwEYavDUXbD6PT8/DcZoDMHnYG/hK4qBn/GJ9mxeMSwRHFbPj
t7kI0vv1SFjwByPuiopjw3mW7to/weUY33HgOQrK6iySbs4yKcd054Rq0w3PBqjRL+LD8WziPpyh
hQqaBcaF+he4spM9HnRMa/DG9vfos6N8aOAHaqBwXcQWel8F7iGH8WJhdrA5X4RW3IkzXSfnS68t
xie60xpzoSM7MYsNg2/4rQpJlz2I0AcWPmUDt32JFY+YoIAcA5w+gId0tBbsKlGrhMOp54JTyUPk
KPWKpTsw8ZUYqGl0vhed/SjDq7+BhPrxsVwfOCSijLLx9yrnQbxXvj231jv6woiyMoEWXr/Ls1Xp
Hxealc8LII5bvZavc1/IcufG2KR9jRphnID1RnlK5iDA0xFZRQ1Xgnss8orPY1XDrtiOPDOERqlT
gUrMavH7V2g8y7uDq9dc+rwlRddKknp8+iw4UUaEcp0HOSaOhk5j81ixADNvDD/7MZpxb+OIuvJg
ziQv6XFO3Yym2srDib4xpveNaTTgeMH3DwbhJURLE6Ye4e6HJZYZ5qZeFjXg3gNuL1fT1v3ylvDC
lAzhw7jkR7g/7D6pToJV6AFc0pBBNj26sMr+DG3cgWurwocdE9a6CFbYx/UBeb8H3UbcJMJI2oj8
yZvd9X9U2EMQcauXNXIsiFWrpQb5DUfrdn4alhY5lSVaM2lEhziu9johOP/Qrkz2fKL7an/ieeyA
WYKj5a0r0qN4Z7ABgQ/FLM4vxJ+KnafP8mWkAEi8/lwCC+lCnubjZU1P3o02J3tqC0kHfURAE4MU
GfUOffos6OjpxHzpeqeKPavdhTr1j7IHvzsG3ZJW8nm92tafBkASkxI91GkqObPUhCObHZG/gTpC
AaW0A8/ikBOn0BPseNveKmJKptvNsl8RR4ypg7iTiYZWK8Ojaw0n/NN/L+AoHDDaiXOw/7rsInma
aTg3/wv9sBrzAJXoeBKtZ43dDor31O98u3DgwYI5eBBoK8FkdZAB5xr/qq+dKa/uJ2l+/bcydjum
ran22XbB4gRHgAGvP1v3CQS0Ft5f7KZBf4URoBdDJOUB6n/1ysFrqUWKHYnm65ZRIXQ1dVlr8V6l
k5XP0sjpMga3Em42fgW1pzRLRO5Cuy83Dp0ZpT6mIlRYHoXlXGRqRNdc342qXJYKUcivtKSmgovT
PKs1Vj/W9RF1n+Y6To1LqO2Q9EnC1E5mGNakfnfYNx9PhfZXLelyZR/Ym1AjDWwxbbT3oMRXvpfe
ZyVV/jois/sQKSgQ7QbBdQd8xput/icTA42sduHzFW16yeW2qCBrA72vXGeg53B7f+keh4zmR4HT
HaM9xU461+RN7ClickmRKB+5L3CQ0D//ztNTcJ/h12D6Gac32IwKPB5EMurcXw8DWLz030w9tfzz
YF+RW1VyI/AB/n+udAklSz/WmV+v8gG2dlDd8qQG9U0RM7V5UKPpnxHzBmI6GNrchGgkgW3s+3ZN
NrXm2aDv6SzOWoSAQDTspW8LlcqVBSOBdDW8Q6E7hcRBLzkBOmwbSd9kVOGxiVC9nsaD5QgF48He
SALAK7qgFcCIqIAE2n+neINcQX8zilYN1l44rkppHIyrA8NnljhGF91M/Rss0igan0zZFPYXYxUT
OI0VlA+5A4R4UTBNM8AQn+NgngpzlHKu8/h9GklcNB17NDbiV6sZdflUgoSN38Ywqba1NjzkfqzZ
rNAv83gC/9ZYCS+yctRpajAhegWTwL3TkoJaNPsnvF65fAK2iVo+rwIPfmtQBtFrRfeLXGixzUrp
TbZxJkSFIV9PDvikX2Qr+vQTNWOKo1vmzROAgEAs0iiD1+V5J2P6VOhdRVOQnEE6H1vMflWCNNJN
fxfilux3Sd7oFepzVaxr0T3hBU2a84au7daVvckMrc/Nji0GbkzKGIHXHw5t/zrwy1jqhHx6t2FM
U1XL6sS86zbRkPevPrw+t8giD84I2rK8GPUonFCndOF7q/r7KRNRbBv9MGDXW3tXMXJwd6A8xRBm
4AZfAO5Lm1z3ArLqvG4WBGvIxH9f7jOFgyIvkkIgc9WqK0XxPVzBWeSZKXz2usi5e8PTsMVenKvZ
fsMNxUVerfwOy9UPtJpRP10hpw5JzTucSPOOS0b0SCevEYlgRgiI8bS22/L5zy92JJZc3wXifLsw
jdEKWw/zZBuC5gCg45AkpMtvn4+o6k4o5IJBnJT8iLg4S0IWSr6NJc2dmdT68J+SY/MsZUAquz2T
wb3xWUOuHLhlYrBOnvvVq3uE4koBvZDi+IFARRDVm14iireoK9oTVR+8WdnLtqwa3+WjHb+a8Eqy
mFefw70oxE2ioV7wHTIqJtkC+9A/jcdNP8TZWCFvD7tiNeOfwF89EztoX+xkkKP5Ml5OjbQlHtRl
RcU2LuD6pyfr3Idru4AWwmcqVMqCV3uCiid21352E1o4L7RwLoHH9NNZPLOT7+h04VczoGn5zf1Z
lQBjZXDpOufHe0Zbo0+tQU0cezq2i9rk9R8ifr0Vsp1dS8qPSjHuZJLcAlgOghxblgGvM9Gyurv3
8FVTHbbawlp5l2x93hQ7BbBp9yLos/ok/foS6QFZi/3DZiQX/tTGe6ISypNplQOtUE0D3essTj7a
Voe9POcDA6hDBzPAghu08OisWPigyEKGuSkRHoRYnLp6524Sy2M7IqhCjqDMNP40ihv/uVxSoQ0/
p5JxRX9tBkFg0rqJOu1j67iZ5nesNs2C1kUf34Qn2Kf4seihhdz0QLrkyeAvLWMm9fPag2qMxEG5
pc13ko/qey6A9o2EaK00OETW+7GSHI7WP2yqsaTCmYYAb25e3wnk/zqPAKELWv8YpcZ38h5K6dN6
id0wX9GVTtifjMjRhhuwu5qSGM+TZbpRZScx36O7rezloEUDu76BvtbecRSQWlRB65eNFfEXgym/
2TBO00V2yBLfCDRV0y4cMviuVdmYRVB78j3/ln3oLmsqQlMWwWNb1dhX9ZpIEWqk4+AwmqZLW/Cz
+D0+pwOp48qpwIz/sAj/64nOk4ohI3YDwH/oWLtIoC/SwyCB7FgEaLflkZk+6pcxEQ6KAimBpai3
RIS/KsCBJz3jq4Wuhxoak6EaS+UIGBrjQGyQaya0UCrOhgwT6AwwY/PLjLx02ylittQ1Fx4Ceyhd
N3bmwusIDCEmuJ80aLVUT3LyRMfsf2Ra5Okavi3NFNg45Ei9pl7Fv0+BjUJZJukjA7fq/N0E7xht
cZRoAwpLv/sLhQwX3XNagYLIj4DxNRIaJnfnttoW2XEoQndEmI+ou1ZzG9NL59sJewRSVYcAmZQT
WzaxCwpcJC6wRd2tnyTo4TtdtZJ0J9gKcpYaSipcm1cKHtWBvaBljqLl8T4s5qhC1jM2o4GKUbPn
8nN1fHjnH0SsP12y6QXWsFOz3Q2XklID19FP5RMktG/fAmssZ8Omm8gtn40nZNDzEvcR7HPRFFY0
d5lzJvb9KOAv6skGO9WDrjGqcUdaW+RvUURYOBmoxsEs74bSVPAhMnhGs+/SyT9/vw3KPc+cUUS0
Iux4juTpIGtC1SDMOOyCIW25tQXtaIyNZzMJQ3k80G3iqYAiBNtMrb/AjQL42OXqeVrbzu42xO5m
k6iXj+HPSxgCp0Hhqs9kzBCKqdFeWTUsThryW5W5FjJyekK+CZwQ1KtAOVxHRjJHUJQ73YVgN6fI
699xzw6b+slICfML/K3+Ge4vt0dzFKEFfxRLn7Vep4u/bRSpp60hf9fkhxWGvkdrmW5PSl9WMaJg
ajBSbfPIQRs/FRXpxwoWMUfCPcl5xWVfygI10IC3WoCpHyrns1gNyytR8r3RAB9byzafVCsZSKCV
Lu9zwCR4tC6zsHc2I6n4cH38t6nJgL956LIo3Z0fA+Zf9pZCjj1SIbwS/+z/jsdci2JPs8JOtmrf
6N0fDDAprqu5md2xIASawebV2brJ5AdPYaW0y46RcpqSKeav7Cl58CSNTHuxpfnX5anQ0sP/tCj+
IriGgmxWNDwY8+3F75TremmPrtEOrqQC98wOuYbh9Xn0h1F9k7KJLw38K89wtuaURYMkEaKBwrEZ
rhIJQ9hp1ue35gUa9UNvDBB3qjFImaksGpSOh8q7NBPpt/0HCV0mRPUJ8tN1rlq09YO0uvFkHhSc
8VqPqE5DaAddruuu95kLJYQ7LkH/xZzxebRmHGv3mj2oaaNCeaNNXSh1JFV9FnEoW7A6k6He84iC
xo57RgcoOK/A7LFqcpXi0Onmuhuh2/Ith4/RlMUc+fD03sGtjOtu3gy1zRzrdd/qGr8UV5gdihDb
AqLlUA0N2JmRjuxmApsOXzgxVUxJVi3mRnnEU3ZTy5Zyfk+syR9nKoYTgZVZMz91P7NQarWvYeol
xR5aScmMqAXQYBfPYQLiENZdZ/cotE69A7B3cvCgKIlXEFzjf2Uk7uYrfZhm+h0HalPfKkUQPDtA
F8lqTO17JDw3XVLjxm4/EugpaORaG7VT1dZXf3sWFWBz1Wo/BgRDyOsDCzCtLoR4awTFCiADQAgv
kotawefh/bsI+4UmEfV683M9gEGJpQHgCD6W9ivggR9HPpwZJBf4ImgBJHlAFLmnLoXb4GL+SqR+
4O7+EZOTA5Pw75Ow5171kpZEer3E3eqAhrtuaGf/LQkNmzNfLafvpAoJDWXH8i8Rcq+mfgiged9K
o7+A5jJHoAUtGCt7nXc73CqNsRWXF08zdv7nyCl6+h3sB1T/hldCHOvfC20BCACm6AvcNkBS6xjw
aSvnpcgV6Lojd9t1hpqi/F2mx0q6RNQG7iYo64r5KMDXJ0YPLOygiQLd+/03M50IRqXSrCHkhh+U
CkqreLxbq6as4ARZ0OXJYhqCsLX02llZ4/VQn84wPMrU3b4d+wAr6TC3NT1OW6IuC2rKqy6LEhYJ
yPSlDyDkateW1XnAFbvZSw1jJRhpCkdKMyNn88hg9n26nD6LrFIGo7lWct2djGdkZRaMo0dsr4U2
IOlRj6gtE4Pq+U6eXFO45hX/H+jK/5JodfNPuIXWH6hK3Do5xoojcct/6puvpBxwmFxjusKeVY3R
/YSwraeczd3og29SVhshjrD9xzQLdKymGwF3GZAK1W7B++mA35R3ymg9GrS0L2KQDuXSly/+PaY/
ATRl9hTTbAO0DCwJx672vA3rGl794xquEAGewp01KlPBazUnDNeYirknZeb+jIPscF1H5XcOnEkP
VxCmjPSU93A0eSKb+iN4/EQG4GidJxQ2oKHZlLy6NFZLtued5HxepHXjNDJqK0IQpooZtntP8Gbw
VLPATGiORKZG6unZoCVytZoEg9rUeb6LpUCskC2MKdQNdrkaaDoSZ+8nKilf+6UoIT+BHVHp6oKx
aAE2Cgo+MPTa7i2X+sxqiTLAvf+vosCrGU5rQyz2/FK1wNtGKrrhGhvxQ/jLytLcvN0oPytRrR53
d+qgobHnGwj2+JjQFZriAIYRnEC2pYdLMPPQK+r8UkB/TTD+cLVpM4QAt3pLiQf6jEGd5Vz7jwdq
z6bhqsxzZ9kUVRPEUM7k93n0qnoXX+Zuc04D+cftUMG9o7SA3bACdEck54b4E/+B352gOhgX2Ani
qy16qBFMLj5usByuNBLkGqaWMuTOEbua5iOS8odcnRSCjaGiTqvmSTjy7NK+4iRwr4JLw82SLWu7
rZTHerxxfDUE2Wc/jhhDmBVUamw3Q9XlHmdFWWunwyG3fKZcPEJw8hQfqNUx6k2iMg1mS0OIzcQP
VInohaxzPS4y00gh6ETWA4Q+nosRZdRpbg7mVRmdGRl2ZQN22V/PQStBRgY7yqwyCdt3yw5Tjzjm
2k+fRT6VNf7yfKEJ3nxVTBRXR+Hs5/zyvjCHHGTx9Dv2I3VBR6Wh7oW7YQRdpBwsN4GzclpIk3kJ
Ts3SOTYEGnxbg4GNJe+ZiEBPU11KFg83bVCZVuZ/yogA3g+7ZuexAYwqDpTMiVDCz+zxsStWxXX5
RVmQtkdxcV+u4KAa2P4jCyFH/xzwnxzU6O1r7ScXZNxWZxh0xZh/bLlOwS9VnXYzIO0oHSnQVU0t
jPYn+Xjqbqbb50g9IfFj/NiRJZMEGyCmmtphfG0s7nxdVNIWU+EPeMnlPxqBxT9kfGlRB/S+5Iyb
e+X6BV1kQkJH7aaXkWhOpSq4yp18s2MGNG/8N8rZOhYjtrh3vC+F6lPdcRCr4u7aSchZW9WF9B5v
qHsT5p1JJmmt/W/HAlBFkB9UNYRAG5aLwvFvdaixFATwrLH551i/tPoOaubqTWjJb/JkIQ3mMLEH
pJV5RtU49EOzvScmhxs2CbNiwaVRIYeOUoy51sSs3bb3QrWxrSQZKWBSaPawUrXHLCugfzQGrZ9+
/pBxWr6ZWkrZ+74bx5WqpIvMsLerej1Bgfn8g2SUkAm1P526znxm4uhAzbGQ+v7vzjjW5Dq8VlHi
+C6c/Sai7fNTwPiLOxMF1dr49b8Z2YyY20kO1ANgDov7wi99WUY1CCcEmTAiTDVK35ge7Fcm5Ll2
XfQnXxJVLPs2dXmOcWDcJxzPUjVw/m6IghgZg04tcD7Ol6yfI/cl8cRtrECZAxu+VmTXaupHqkxs
wUFlWXmjxBke/warHOcz83qX5748RBehwEy4vGighJwbwQAqBJNfBsnz4uRdnxcQmHcKUjbY/gqB
MkQAd4931HSemmLB7qSdTOsKUpAqvt7qqSdLS8D8/azDZaFxDxMMKWDXqCcHsJiXc/Ydhsn4lzqE
9fj4pomrKhkrw8Y53GnloM3K51i5vPXlDDssOOZTHcF+APJXSUckxSe5rVVVYRR485abiT8Mwa+2
g1k+PgocaC2uG1EU88L7w0H+pAmCofiFlHsR7Dfmptte5zUW1RD9xiA0SvqCy6k8zU0xorEvr/V8
Wy+H34SOZEih5J1hkd26u9Xa59gEmDyD5M3slDfhpnJwDMD838KUmnl+vyMo4+AwsYwloRGOZE0J
jo7TMxNB3uPhjhXGG3pI4D7Nq/1ft0u48R0mWs9FWn+3E8HVqaq5ecgFQ4Ecmn09yfm+OUIx/3XP
TGu0ce9yK9R5zpQDEndEosNm6U/jrSNLMe/k1+MJp+VqD5KQGGotQJC5vyOu9v2xGx7eEoxFCv87
P81HBzNYywUtdiHCHlgeuX9XBB6A7YkAcMKZ0Dr452K77tGzmgDlk8lss0r4l1OphxWTKC3Vlz/3
mDQe6ciSk0Lt/haOeF+Qfc/PTt3gH3nbNFfJfFKqiL04ioHT0u6LZZvdmYlfR3+D/j9wlehop+d1
zG5K/eYr2juO3yrVePIFG1D/M1GZsu5v1R874OKig/Tz1GQY+VRoUkouVwYmR2U8xsPtHi8rXFsU
Ys8gyK85kOeOfd218DbMrhA7b66qMtg59ZtHt5mWNFhARVC31j7dEeAOfuHtDpmM1DKj3s3TNc5t
x8LH/nTUO9mSKhvP/QJxm4OgfyfO2CQ5WdTA12kwaNXnhy+mVMA0+t0E2HCTSdxa4cZaw33GoBNx
P3Gv0aknxgXijhEx88RcxTjaZBXF7IpAds5i7/yL2meQKvnCKSzim+LGyIcDRqH2oRerOHALLhqF
dJ/58DwRIApONv6DwugRWOCPtd/zPbdmywVAU9VdX0dKyPlkqt2KAA9Ma5gHWTCEdhG2bzb1U4YO
5o63WAe+86AC3xhdfeYkDwQJdikpZb3FexCQSjyMrzPmechS2I5N8YhHqazxPAYyFF72SNfts/G0
/JPF62fmC11pEe3Omk1dcLlE4MvPaZ4AUoZM1f/+iWly74wqaEubqBEj60LqYsKo2arYh9ftNUs0
VInP5QQ71c7iNOviZgakaW9FenmrGAkhG57dDds3FoXac6ND1yIbRS5aSOUBXrxcBCd3fIVKP96h
sTLWsB8oGpl7MCkjBH+kJWjQKVU8zV/0nxgcMvrE8n33HVOlNPYQQBMSXJWvSb344VY/9iDdyZmr
6cs2EQuQjdt8FpMjhdNmaL2grbU3+ozZHWdC3kbUikFmuYttlTPm49rEelAVOPhueBhZhK/IvIUJ
LgHq0td8rikDZ4kZ261of/dzuF6D1PwHcYTllU2JHvKjPPl7ctI4t4z1lcoowHKtbZZMp+y48spK
bHUdhfCq6IVtqj9lISFjpiMSN58uB4AEPIh4vHk5R8TUZ+Sak5OMTh5LBmQD91gMxh38RuTzIIa3
M/8C6Dj2LnCAmE/NKe2x8raaRdyP6VWjt7BekaKzz0eyljvICRyAzpAQQW9tc7PGi9dZfAzf/nNs
tySsrssUsXHzwvhk7wgSpZ1bkFpxL1AbtDEPTg/uYaLOKhPR8LmFfe66GRXd4WbM8+yQuuwrgTCl
RM2s09Bgv95zEFNXU8SMselyNrnyxu5EJYOrIyVIE4wHgPO/tj97b5UUC6aEiaWhnOLmqRZB+Zbh
Bv50dC3J+3SH8U98B4QgROxZc6u77J7g6TvqBVu6hJhMCInrhKyJrqBslYuWuEoBjmhoXYDmDNzj
v1x3rvKPhMtKrXRcQoZNFf9aWL8eekDHM34U80FyJ82W+s0wlrZ+GR3iE4mNiD40lsG3hIqc2Ekl
/R5TlTyeW1OfupGwUzCu/RQjaYjlPJVVWfoNhesRbv/mVGq0GCko+rAlkS57gj8lVtG1PQay9eO7
kPF/3Yr0zAWuPZhTULAq6OfVx+/w5FBNl9XbEnJhqCS4AppTqo+HeQL13uKJSl9AYDEcdiaKXoAl
FBa/MHdJdzyboM8yx8LJnpcBvLpIZVSDkHO89zaupFh4PbpeEYBNYDaZYz9i0WAJGxp1Y9iOhg3k
J9KkVA5+H24NHyTrv7K5xlrMHUjhcm7jgyhh+m+s74y6ErfBiYhgAAOyOnbuwBgqNftS4cWswPOX
7WqyzR9QR4M88ChMG1PFZu4YZFANV+dvACQEPfBqhVIlTSmHIBI0fwEyKci3AF0oM1pPHr0yD17Z
NXFcdaykQMRfGkwKy4L79PJTfDnSUKVTJAYrnT6Aj/bNRyh8jGsh5ANFACRNexxzH5nhlgONSUpY
NH5nY5w2t7oDNiCdEpAM1Xh3yjOZOSdQO+q5zILpjSUx9okeylu5S12YyhXtVfiNRMxUzWP3bvch
0mRhVxJ2qrugBgOIIcWp2NZRQZbPsJ86r1EsW/T16CaDdaN1Cm+99w/T5KRGUXoY2fzH7Fyx0ISz
bNL4pBRKsg9Dq55YROyQ4KYdgJxj5C5E+oamEm4jzZhkNNirdZpw+Z6xcmt3DSiy8M1dMYvH7/bz
Qo3r6otJEUVXW2cujr7ES8tFjOmytFH3qBKkuonshf4/HPv6KfH2jHVDm1DxSCsJI5ecxL/cIJDG
ToP0ELUIUJOPT8RRnCr5stlKvxkf704h8dud0JvkZgeavZFzlMAonPleYDA/hbdCNp+Gg0sQVSMa
PfxPmfsQ3LONW6mRipRRp5uTxK0XTAKDf9n5EqxWzkhlRirNkrgiYlOEe8XM8QTeVpeMVshDGkMu
jfWOxoLNCVRgXZMl32COjAwnOnfKZxXC+oOuviAOk/KY7ys0ou19fzutZjof6goLdugfQ4JO+tgk
VHuWiTglHSG/1SjlNZRurR8HiF5XLX/G4vQW6xUkWm6Mx6rEyjJ2M6nvc5imr1E9DFh/puw5RSwS
wziOaGWuqOk2Wt0kj+8RsMDoHY+4BG9JGILXfArxNFIbXLGavLZbtvO4OkUMubHz1dunJH4weiVt
mHsDLnlpGOC8R+rxCP3D2PWEgpdNyj6lmIXPa6YFKveI7wH2yyd3IOrSRE+xg5dWzs1WFLrwDFW4
zoTIzasxblPA/8OOhSLVtABcqwr/piBXeAhpuKIQikZjDSijHdy7QqKYDy6igu/5K+3rdberEsa/
YQ/NN1Du/yLYfxiqI/wWFTIIDzFyE5xfI7Wo2Spgo+J6jC1hfR8lVRmSolmp1v+F3zmmDZFAFTU0
kQcVdCdTOrrp+cC4nAaV/aj0tHqDOTo7u7m4radq0jjXQfcfvoKGdHaGXWzwvkmrRnbDLovgJH58
ybV6vmHuIGMiBmQ+j3bf+nqqcJvW65Rl3LkXvwTCRtFty0B3gueFqHiZHs89D1VF8TskTDWfWTnR
ESAkxvb0NB5fmY+UUw3n72yVSGG35qnps+MPrM+XoCRHMBUVddrikgCPl9i6mKNgluBV24m7fNIv
pMLfu7zAlQhr5/phRC4fuoRBBGPcja46LUDczY8Q2taBMeAFE9eORjsMMJqcDuT0HJ0wSntbo+9o
PD4DeGmpZddZ5+Pbl4dcjDh5oMZnowzWYX1Ms7v9QqtRKfjO4dsZQiWeVZ89QhMAGsX4uOI10LDH
5EPO32+GZn2iDuY+naLgUuODgmeTJqlorTBktqC2MTvVnHT+DZEdL8BATXyxDG1makC1OsDb6wVK
nDC+fGCGuhRfcbCtQT1rMVxDhp+WT+n9IiUVd5wcpBcuMPoViwYNISn7mQI+s6VqUE0jvrylX5F7
5NnoLt1PTSlFiiqV7OguESUvmCqfIj4G+nSRF8/tzWf4oAQzdgQwvyyIjcxGVidtHkqeU6jhPnR4
pnvvLaig6DFqL46DPL6IiPACiaiK3Ask7zKzynIcFCiWPJ8vzddsK4kDCBhK7EXHqKVoKp6RCDD6
tFTnc4UKHeB8hGxdgLbhJZSmJVRbT3JPH52VU+dnCiiOMaIhEfJl+D6bN478FgXH6nC29JjxFpWr
0xbVb1zunpaxG73nHwEoBkojoW4mA1lOMntQwlU3iP83bwwqn92TSLljj3xHZubeUEZD/r6ffco1
JUsFi+G8aLfEdnt99HDhhcU3rLGWArpH3QOArjoNU2MfSx7h/mh8iWh4gg5I5TMF5bKRNrYCqYob
pw6G50hDQezdHjbTHPWjBc67o6fv9aJadF8udo6YNSGmoTQYUGarCaxMXvIANH0HNQCLEt9paIoc
ip+h8pJDdsZRKia82932oUMR940QIzfdb5a3gDgnhZvFH6UiVfX9bIErPzfaRtNnHRKrx1/1E+7o
7sN8wt5f0pWEZGp4ps6QdkuA0owKSEGqpJqgUW6SiUePcwLoyTY7LagYhIsd9EtbNv70UIDVixCQ
/Xf6JMDiQapYgx8wjd0uVXheaOC55EylV3aixSj/6GDwpu2ivpJI7oYDvCR7YxknD1MPo5oGGeKe
LPa9Z2w45/qaH6ZLCtAs/J4eM+W1WoDtgIrQPSE0fQyzfA422avtcXJ5i2sEmho3FdfzC7NBwshD
/35mlTUjf44FtF2Fmm9K+8TZdP75NMRbf3HdZpEkIy0bNSd3E6zRhRM6mZR0i6gKOV9HjcSfPMxy
mehU3OqjOx491C0SP1JBb3REadF7kwyf6LC++c8xrUUU+A81eZaNbcyXkpL/VpPxJS1MueWcOtWP
xwXmxr0GtUWwkTbxlQub8Q2Nsf1UDFmZkjBpcDX+qMULliNOZhtmwZ5WmwzV+TqBQi1oWPmRIbnx
QmHjqx8wGb7zipxiHxVb38ComhAtqxwju/0jOOX9ybecwsg/CCnddU3MO+ZVUm3krxw5f8+p3yms
16kG6xANuoLxQQ8K4OdqaeG8WSd5537/9Aow2rBfrbZ2P0J7+PE9lj4SLRkq4A9Yv4qX1QPgT0XN
XT4TTiGxqzmYfDmShnZB7UKDpacgrIBASMSnuVXHr1MOzBfc4BWTHaHFla3QwsJzyfv4xrU5BfEg
EPFXbHxbC3yL7q21Zkf+mt8yd3Ih0yNWeVqPmuuDrfbfEwGHBk0IHANpEqr5BA0e78PJg9CsLMih
9l21clVjnyLl9VcfC+luSJSDDc94fdRD90jnbeRfIFdfprO0zIv6WGwSvSsGUoD3KQ98DlNYi3k6
O1zGa36yOyTgh1kHfVD3KDPLCtrnrmBBBVzOpe7saYj16NGUSxqxgEGncvI8o7fVIzm26YLEGzPK
ykhgGVleP9LiBRMggu+zFfLDoPZQouSD61B7FELjIZHQc/2I2uUPsmMA65GJpk+Gaoj5g9zjH00F
Qk6Xi53vC3bLH8wAivJoRZojoK6+YdsXrC2nz9c3jEOsgizn9qix0EbqoBsiWlw8Q8P6UTJgTCuW
7XlHcVVkdYmUy+IVEAmC82XthYpC/8WxIRGwb2H45wIo7bVYRTOZJClblCAr8czwn6+rk7igb3d7
NvIZXy7AYqkgFOnSN/AOU1zILx2KeQQGpfd5MrM3JMXlpwW80KXhQFIo2jox3GO2HQt26hLskPVV
g88eHdR4JpOMPrE9c6rN4CRTMwT0IQvK7wG46Umg9az/F0eWGhosan7KwdEQf1XbrWnaMAbW+Dea
c7fl4MPcQGoZbV0h3UtCYfyVwETAcBUYdY4TLM4GPwV+WEgm4zZvqWWSDv7GhjSmUFGFjlENge76
4Q7rT9w/VU4HR2JdEljqaz/PtjfQe+fen9oQnTm7WrvHYSCFgLV6Udo5luacGhAQoqpOXxpwKixy
cJMdZkGENfKssUPpwg1wZAkWf5fQwfB6YSaMCvYtINsItdPFKF2CryX59NrSdjeyPuSWtIhONMAR
LAcQrYwDtkpTI3BAGtLi6aIaOGuw+5a86RZOriQGm1trhhYMLih4FzdSESOvM3bG7hT5Zzr3zEQ6
s1lCNZ3NJdzPZR2/sJpNqQa4AGOI2UpkHbSVvJ+iW3lvFzNwPoohYtf/6xkqWMn1zLm6ZMTIfWrQ
zecdZb1rIWrKtQQwyEWbJiZTsibt1pr+KQgM/+Sw+3Hk1rfD7GLE3r/7EUe4P5wND2x+m2tQ9DJn
w8V2jUPKKJF/TikYM5EZif7l9/fqDmhBWUsVvmjbTfQ9wta6Lu+6U6cn9Z3HghRKfVXoH75fTLzu
qjd0IsCq2SHyS0/IzjYxh3Chgq2sQ64RQ5mbnPZ/oSnJoeul2KlLkIfXg0+5Qn5z/H6xGsx0hD6R
Z1mettBdEX79JcfGEzjvYF11TIUgjSWxcRipLT1Y6/JJqJUf2LZATqeDw8IipCv0EL0DZavStzre
WuPqHwpnqgTXBbYKaCBpZ0Eu9JHZPwWcO8Mo46HW2CdCoMwT+wd/GxOoNs4F6IfUg0SnZXZUq3ul
mx61eYFHGg41XCOzv72refBJf9EYj1od6ZRnRQ0bRHhruJCRmysDFins2h/GKX6clyWKF2RFPt+w
PwcQEldKmcTLddvYGlIMIvKy/TXQ6fMYLCt0TZOPFeuCgjv8sPmp6EOtx8up97Z5vS9oROxkBgBc
Ja8e72PMjkeQXbTZEHSHfMBylIpee2n8LT3kEE8KjONuq3s60lWwkhXWed+sv0RasKQ9ZTEaIl/S
KJrRpQ6PQIJXHVuGcZ5S5L+Fk0XZKS8dZEoX8fnOS9Ecc6oIVSXVxw4bWWfG5c3Tk5TUTGYdgHOh
jXHqoppZTq9l7GPPawxMk8BuXjEzfgjmkeqbOp3q0AdCulWEOQbve1KCf8t1A9VLWAhycp76nJHz
0gXmMFydXetSc88HUEzw6SE1umO7zNrXbVwiToqoIiwzLz8VMosKPoza2plu7S6DpYLyCiXPbEr7
ZKkUJtKx6/pgU8BBz8W0GpE2THGmlOT1aT32YJJMl5/ugA76X2ChYHJqhw7pCM6XKH6GInC2JxPA
cSOi+etoHwq9uCrBKN/8aRzEYCLy5iplo3lwyhYkkmHixMX3Dt+cO3vrcQ2A801o6UG2PiLvQjzN
8SVvIGr7fc+5gzLbPt4sVZVKf4ntZ9WyiSsfuzmySZYqFlqXtfOUioJyq+FFaqvKeI+6SIROO+vJ
Mo9q7kkeHFASZWhaammqiBtk6nBHlNVXrL789+6jgPOsLGytcPpYkGIrsOPKzY63HuCutOHVcsr6
tWcyBiR/I0ShHx0m2l6vFkLHmuHZjdeUFQ6a5P1Es0EEmteP25jOSieqQQ1xIntDDWebwKQ6sdpc
GvFG0i6wWG56w1vrjDqhfklaHXt+ReE9FHzDw0l3NeyH8ww4fobKYH8C7a7A4uDJopVlw6YkaOOa
SOZEKVyuN4hshkzoGfwuX0eWV0SEe6b8HqruoL1I2R39UeB4AigAr9tvQo0863FvP9iouXrr58kJ
BG4wVn5OitkUwZq9mrAUkBb9gRkZ79rOtpRkLuH8XSv0naFWr7YP/vWHeliBxWJZSlePfuZqBwoW
K411nAmu4K0YR85oLeJ6MRJAAhBkbgFB/TGGmli6whqVzqVcesE57EXwuT3c6LXqdRpftdg4offv
xlXsieKaK6LQgVX1rDaQTbvkt1w0thFqG/1rGGDaSaW5hbrKOtdAkDRqZzKgacn1VQSo26U6moid
yZol6jvEYlpnGQALN5UkxVbhvKBCiZNsUVEutx1qqZf75wUfS9jti7P+ZhHflkCb1lqvkxzMcGxC
QNcrry+HvzUe6ui/F59KldAA11t51+Sa74GUJ5UpBDC4r2I1+SOEWlg6q6aJfy5e6IudiRM3C5Ep
27ZzJVL5Xln0B2nBcERyOPc/zspbpA7vcbPkoIKwH7TTBDrbbd7kA2b/ee7SX55WsYdsplEbLawe
zrZTAOTt/wy2xgcwPgOTcCVArUjOmFBg3EBkH8QQ6D3BP7OpCZkQWlz8iA76D7MRP+TbSeVkqnVL
MvxKvQkBZT4x8gmkhnHAP8kUqzB8UDCSAotV3H47oKi0r1Rvp0sbUuE9u3z0MffYHj0bbt9+RoLL
/fJcLMuq6SPSroIk+z9VyfFxWomIWOq6CXtOLSVXf2ZYdb9YNatcAxtO+Kj8LRfHiS3JxDdvl4tR
lnJiCm+d3tM4lIv71IpPzQtPBQzkww8wc6N4IPlYq1V/t4EQ2djgl8BbIQdomGmMIH2vQkV0Wmt6
ZUloI/99rJB9HvLdMaxXF/tPTp4sWdi64lxTox97Fg+wUloqOda+KJmgyzBKt3vFMWJwpJCZQx2Y
MsqLUiXi0hOojHVbWV5sxcVLC7YCein4wU4BbP9w+wrWi1uJCMbPAKyAejN8J7fY/h0zLzYAoq1Y
D88Nhv9+s++Onx+A6rV1rh9PHbHTvryv/qhIVGLStZg67D1QqmUWwLEIezIkxUHta0Su1aaDaEY6
MW3bnr7dO75X1prODulDNLSHJFg7GC0KsI1GHZMUCV9t4/QFVFz1nmaZxV8v0mK9XDH4kl/ani8g
3uFedbeC+B6K2XMokgUAqLJe5hiFYHXAtRvXLh3a9uswxxehLo98tgqzXHRXLsA6FRheAfN9Exlf
CRnGjFQxp32eGfnWsIE4WN0Nvy7OcaHhfEBiiIFk5spxc+x2HUTkC7mDYXq+xORF8WjWkKwogO8i
rdxcj3zCwSke5Zhd6FUoHdSxVDGX8Ctc53DirmsZAh8vbBTFCF6fVEAGrHxMpYjjsEb99DT2vkuy
7uFPydftkXG22/CxjHAktA3NUTriIJnevyOiCBATWCei42J7zP5IHKQrYPowkFsnu9h1A9j0fFGU
mouPH9b4i7m+0ghbhw3Y2LwnyNTNN2o5fBIPyuaa8GHTMckpap7UmoSfBFQOVnAHxGtAc7s6p+wl
WUhirEao9HcmZOYDj0k9VmCZ0xHkVHdEPFaHOCbIn5BNyDIHhYr/bxZ63q+Os+/WDJ75CV6P9t7p
yBiStW/OECJ4kKfQ7uZPBdfd8romyiu8hfexbUfVBH9jcYhTOwUKECrQnS3Wg0J9oD+dQIAHPyVO
qVQHNzRGdsVmjOvKU0oC098F5TBjllyh8isPlBlnR5+RJnEwThn1orwXoh71+nq1KzpCwMpai1Ux
cwwpfVbzlEJpQHMUoDWrr8A2RWdexzk9cmx9BJe4m/YK8t3pGOmkOuOjKliOCvRH6/zkJ3qKOHGF
cqWFyR2ndY6NjvvE9gZxRosVjaKh1zzRnAH43xDjMHOhIT+BLifLrE6OCDoaR59s+V7mQ9bXVpv+
kZuDAG/iRuSb9SEE1HIie/kSjmOsscLSEfYhV+ldZchhdUahCizibdiRYTlWuXkacyGpc0Ocv8mk
nA7Gvnq/RJLIYC87d/v5bpVfLXweRylxUXYo/Ym81Lm2TBtqyaQfuyxBflLifoemRtzyF/k/qGbn
uEzEEyuNopAG0ICakrXkqHUXai2yi8a4Kc9ckencptVczw2vXB+8OCptynKRyZQb5j7obz54aPPm
Gtyk3JfB7mVQBzVKUAX8w/jDMkKwyTs+JwKNf6B8vdydE4hbTEI914xvvusyUjmEh6C8UtsL35KB
jgySJcJYKaLf+iwyPO3oCH5m7IaVPn8jdEt1R6xW4K9aaIxtf8E2HnPDXRE1etPVu+D3EqJ7m4Du
Qou2Yk4O+z/Tr9E0crwbdcV0E+gQlGmu/F80pxYkx9Q4ZbtPRaL4FNQsXjXoFqhNLQ1+JQtq2ZGo
U32W2TOzsndp+NXZcc1/bVwspwjhfCqthEk8IbZIGKkdWiXD+VbUT3CN5CXs/6y6CsIL+omGCPHv
B2SelWFJaU0E+vpmD0F4ArUi2SmEl0j624ZraO9FBCS4AfQlEB9MeheVtNvKwPVYz+igK0iqtdXo
TEEAr/y46d1ZiFsWkWu/Mw3h0ldmSZ+OnLXaytJ9VwyrmC5hbxX2iGeHvCDrt8klxLgkLmhxbEKr
vgmpnxEMKq/0XeDpH4ITMIWMVqn8p5jTgl6cEoeqn6NSJ1AMtJAbrzzhAy6pIjca2WRfNSOE5/ur
bKLSfYB1OEz30A8XZpHGwh63rf2a3yUYG8GdXE+YZBWs+eTg9lTpKS2e2h9hQ+8o9L4LRT8gqiGw
J8qNKVt/kHv96zMM3tqyzzvb5KLhLmwxReWbcteF5l8p3iC0ZmeIaoj2LXmPMe4rVkeLgDSDRsiq
kEzaWEdaM3qvH7dGyvtaN1e4w3FzQbDHc5AV7t6ZSWoP9GHdeBdnUQ9k+bt6NNQi+FYUwAfHhh2T
/sS8k2tT1WZh03kvdCcdzVs5Bs0BG9qoGwWrWoNBoCAzp0JspZUkWhs73WBo2feQ4jqD0Wzl63QT
y4/dSAdUASAWPC/xOJuIkZ3DFSbH7xlHV8t2VBQFcIhMGPxWQKYbk3Xy5y8w2aLP4NkOUat50rfn
TBLrC/w35BKc5aSDmSzBzKzHU4IHhegqTznG9tO3KoG1PhvGQMuA4KEG/3ZwWLrMmjoBBT07CaGe
nSVCZdzEehSA57Wgdl9TQHC4rt+ByjKScjmJxcBuv7OVoq/0LHQKrGnyEmnioPVKtCdTzx+EQYM4
xxIKoRyZI7o+uO4Hr0B6TEIFsrj0yKNCWj5IKZEFtAa28pfj3nRxw4hKBQdXxKmMivX8zYphU7qH
DH5SsTHbEdbshcefwJtgvR00Ip3PWEp2grovjalyyDRsiCsiAI724qyt77+cznP6VfgRdnY2ewD9
EtBZfKG51L7kuSt9nNxCPjb2ob5PciYhr33Vav6JWhGkeBzWAmX2mVOvrBK3UZ2K2//byqPSCyRB
haKZVE7RANPT4FLOODmhNgAjgOYY1uxVVAGsvl2Aji3QGHbyjm6pLGWG2ivsYyqpKqz/rsWs9OWq
wf2iVy6dhaUyRT3pGiNBvehaffqOFuesKiu1Ticza+PXjnri25bDZsu9VSV9zii21178P3xoMYoW
Mkoc7DItlWKLc1ZO3K0oZhUqzYcseLhahd8yhKjnv1ab/oQAJdC6Pw3MlHBP7YP0/XNUETg/9PyM
OA0MBgRp5U2fenK6GcY5+JdwAxu8Su1o20rWwlHv0DW0qWc0dhmZYnjHCNvsixdSTbKXPCG589is
Zqp7XPUSDvIcP/mZZgLJ2b5xL0J9YgPM/sEzcZoP75UxzHUGKKNCHrkFlhTVFb7evTL/nEJrYODW
SfAHqCaWQAawROP9FtxEGH+m5o7DXtIapjggH7kxVu+QCXWPPaYzyxx3AwD43SSwWtsX3bX1wZTx
g1HoUhtlnze64qqYayGPdx2SI8y9ox2KF0Nxz/dYqa9PTASfEAhWj3K4BA8jJpMwJmzxvfiJC1LM
IVri2D+WnUJ4UeManAOWVwPbZTC5RlbambMozm5Oy0JcQPzcUnHrIGUP8ttWHUQRNPXtmpOBJAfz
H3+3mrqezBeFuL05p9emRu0OHCGpoy38KR5oGm1/HdRYKXsKyF/yNQpJvBeybKHcafVvhPwQCEMw
qox4AIZrde1WAN8I/Fpw7ERs/TABmtk9yetP5YVYuXN0CAisBEA9KZqps5QeufhhlNDLavRNTG4J
bA02WDw2d+qBmmo+SxgMlz+b4TnyIVg3ITdi8H23OyPZA8q24r3t1stszEK3vxAYhuHd9T0F7HKH
pJFk4mutlOqemC/Q4EWSOD8RyfnYRPTBiAwKnwcVA1ZGm+Q8Thax72d3YE6Kbkr7bolkiOY26Ryo
R0MzP+PUYDVtj2UtL4kGfh7yFpPoDZwLLwlmoDrhkedi2PK3sEnr1cTFXyxV8KSEk6PMSgYHVvcI
GIpLX8KH1kn5m+uixHH+WlkMy5DfC/G2RJ9fF7rPHIPFBCycIo6fGQ3bZkEl4DcxS74c0KQBVcmX
l+qQngiTUbNeC++c7LbGN204GlRotyQ+s/pBS6rNZ0zIq3unbLZGKFNFo+RShll8tBcmaCutpL0n
KyYGsRwuBlLJ7D8VExfDijVsTT9Dw/9+MjTlgx/XP4/C9xyBtvr+Xc1n5WFwqSPg0f9Tg3iN8IPV
w5i2ngXHSpJLP2w2W2FVslYOTmRvyDLqXwhD4GMowD+q8FFIX91Q0xlv5iIf0/hEfoM+fk7bgyv1
ZZvuGbniKnTdGnBA0SUF7cwsExo9bwWkOz3Tn9OBiZEUTWHbvya5B3qo8XmFTsGu0xLcFK/w5CIH
YRT3eYO9FdCccd8nMshaXN2Zk7ojqugunA5QORKzWeoUMXA65B7dyxrYC/QTmBYy1IpEZIHILtJi
jl0fog7Rrd8uZSZMoWvTQr5N86cmKfSdpOAsHMxk4Uisfxv8L2e7lBCMjzMxVDDRwTLgoANdr9gH
gACovTXNUT3xj7EhZL+I4QsGX1w4wFkCLAeFrYldj/apqTWEu4Npv5tmkwQTRDA5O7Rukp+WOnsd
CusvHnibi0ndzoWMqPA7umur7XwXUzYtBuZmrhu2KfiHsAbtELl0/hY8xnfEfxc8HAMX6q+9Ybyr
WAADFQ7WT82jgoVxH7Yp+1W20oyJbbrOgt9npxRLpCwYyt9UM8bNBL2l8Wtu90jLjd3gmetm9F0g
m4XEv5jWZG7j+ytLG/CPkY15xGTGZstTrxSxDV7rdCzoqMdfELcx6cgH6Bc6HvV0pac5fJAEqtoR
YOdUsytLowtSwM1aSLPmXN04lpnB8rZDa0aG95xCfTu7an8emmnJC16CsKh/LFABrE3RMwJjhwQ9
t9Km8AScdkt2RKdilQG3FyBnazOq8Trd4mOdoxHLmeXBH6C9zGXucuRe3sIfdRdksCdTx9YB6JRw
3tGP6zmqHIYRAueJ1i+OwRdqsNYZ79jwDYbnAfiAkLf398SWIDjVfkEp7nOljWYdLA69PIf6YrFd
AwMsNNl+fupvDuS2cNdj+F+m9VqwJzXiTGL0wSxP4ZSzlpqjrJXuFJEvBxh4u4obqB7reOhIFY91
NF5S3IbP1VKKyurvS07F3tZEWPpN4OtPEat2hdh5APW7taOH4hDFteNpx+CtlZdnabeD9Q8o3mS/
ceOFft490HpVo26o9A3GicjS1z1DmwLbnTeV7WczpifFP7i6lRooWWtLj7/+8VopwF8t5EjjZ2I8
9+VQnF9LaU6VweD+lf+fidSnUNnCBztO4bb9HenLHQAdM1n8ObxkZCFSXWbaYS4p6xG67W5efO0c
2uNq7LHPKTQe3TT1D2QmWdsyPc6SgAPUKpG7bCm314+DZps7K2tidjCSXNi98hVKm2OXt6p/jMOL
EbGGyyhAj6vukEJhMoHWVqGzhGfL9c33/OWemXt3qptYqKfxylEyxAsfDFCNzfAPQRJlmprZo6m4
pplBo9RkuAE0MaFKG+PhoUZYFmaP2HjsM2sjMj0DGoTy8guk4cz8TPLkjrTr9ETCdCzJ1hwsT3PF
rfPW/SuZgNaxfGH0ithT7XyN0fX1lWKYqiTGHhZQ+MuiX9p7Z9tz2TGGLfXeqoahsedE0MKVEMGc
AeN2XNcOmjy04H9FDT7fAHAh7pUuN3cBXyj76TdMAFZ/QqaqEZ9C/GoDToq2MKbOBy98xCrordEA
KHoWjDBZtoNvpBJje4yD975lZvrIVIqNV+hmslj51BMTj4PFQ8h9tXJ1See3pmPTvJv2Dx8Yrbc+
2kVcE6pfcRMEhbRvQHvkSBL40WabkY8WVlhhX4hNQowDrYBZ0Fjrkc9g6iXcQOJkZ7E18j0YXllW
I1J6eMX3QjcdKbiJIEWGRegEqvSIcxwBy5ofVyQwxrBQLMYwKucR18KX9w7cMDcy3vLLoYi+/82M
/kj1e8ah/nWEQAYnra4864H6VMycB1aZRwAcuaNjp4kADr/izhTdtn4dfkQnHTJUmpz4QloSZgGp
kBKBXETaphnZndMAHvR+qAZ20ybHu/Jhk+7PsMsvFwQM2uFH08w1ng6ijnYWtKaflIuMyosz4wFL
Ckp8QBMrLPweY7k+cqpURPVhtlhVFVc7ALIkRtHNpxbpZ4kMHNpJ07KVxvztKXK5hwLlnUxIrQOk
k2kYTPJDx+TWpsbfKg96PN2K1XcBX9Fh6oDcMqpJRiqrZ1SXfX9O3bZrnzxmucBOGVuuhPzcBi43
1niUIPzcqANjg1wDCcb0UhV4CC5OAvoltEpdeem1vI4wwvFAdmxsJ+S25Rv7UEuPfWX6CaEOpd0B
HU85JaWyOYacw73NqlBm1XtW4OHze0am4t9F2z0S14bIjw1j8ad6iPFrWEYWufw7teAqt8Us/SN8
IbYxRVy4qU6GztdfHcrQuayY9Tin5h5M9comR/0ixrTyRSWXy6PZ+SR2APUDc7OpZ5kGa/dqLeRi
+xEjeus/vj0EgwDU4SCSMBPkgTULcLhQ45kkWhjQpnRI2+V5x0jfe7Q7nXb9GcWizFvtOVw83GFw
69Z0siku2tTJiXMEWGMQpmMayiuY3khKjJtvrJ9+HJBuVYTBxQFwbKcKLrlhsUexUYVs2dtekbtr
8WMyPUoOPbSeWv109xsTtebtWZggHdwB4Z2LCHY9A9QwsYyvK948gc8RcYMH90ddWRqob4SnIhlE
piE6VBjYU4Zkm61x43dbLusEfv64aHAjneEZH+O4eFZaK6Ls9/e6FvoT2dXbV2ccCTAwdVIGi9lr
vg3M1vci8T9EQbiOx2A6cvlWG3eOrmOIcXFfK81ULR4lT6wb+bU9cWCvpWAvk77B620j2/tTHck7
halycorRtZHuKCN8GlljFPsG/i1rfZgDRU9nnowRGx4kFT7uE7HZZMDKEBqolfnGA7RsGh5w2uo/
PDavK3g+K/8JhMMY2b0WbOpc2r4dOAEwNL2Xm6MSs6pWJFDZJYMGgWHguGimtzlnPWpuuCv9a1Ru
P/HZRtqIVF1eRT/ui4sxSP6a4ycrBw0zmFzTEwhbtM6tgrzfqBAcT1ickUk0JaNu3f3icZIB99mX
C6G9uaMPok3csIN2OvrxAM3MrJrJiKQwSfwmYoHn5IyhiRBhkzyVp2ztZplzrW+L/vxnWnFZtnlN
vPcMptlmgaX+2MY3mCcMBnWN348htKLJJTlt9VsH/Uu1cSfwV2BDEtEudtfrwUwCrsbyEx7PA3NI
FvYsNLrhptyjU6HgY+Bs4PGlJElBF8/omugBspyxB7bGPqcYcgT4HuXaM3CWfCC99Uli4AJUBf3U
YrJLAxzQLKGfkK8nNdGfAanoYeICFb6lUEmgbXD3ZbSUl6vOyUD4q2fNz+zUROzZX4bxtjshxAZv
oelTdh7hlKiTZA+Zt+oyCMX4Smo6um9lV/nkPmZYug8qJJKMiTzYqzbWIE38hN35mR9Lavt+yop/
+a7koVg1Jiq0wFegwJgdKMkY0QVbpOiw+HvRyMy4kFRFlaqF6xJeSTFDoB7EDFL0/G8OmFgiLScS
Qb5M5nVNcKsmDieSSWCDXtuuqwl7OYxC3+Q4fNBKFZWwC2fGi/u+9ePUQccr8cVZOJdsk/hPaGga
VQs299xV0MjsI9rqywb3gXUtmU6U6gmC3VFKxOXF/p56ScACMT4tshBek4YxIQTvh+/JjCg/wK7t
ZTrFpMYzW0L7Bunh+4h4Ok0bzt3VQDVzqxqrLklY0U16esJx+7bOO91v48DfeJ+gB7+192M9M4bp
YcHAxHRYOt9PlJmRHg2biaGFaYvsXB8d+HuAzrF7M8ViNbBFRGjDFmht7Du/A/cyixQqwKkrVB3a
M4hYrs+X0wUS33X3DVvTF71jGkWcYFuqS8fROw+POXptTWUnO/FborwKVGucdOyW9yRt6cZDGpWh
A8wno3cQkZbT/3ZRgPhlTD/oktXpgzkMdceulxKXFnG6MTkaaQuX0RahX+3dG9mTKyjvwNpKYVfg
gWUBHaIaNbE66qFaEaOq6MNl7+8Q8BgaDHjHwBaBHdEzsaQA2ATSAma/rTsZ64L9FdQPzROyiSpY
TyOieRvYRLoVoksFD2fhkIc9Pm/mSw0ii/w1bQFU8GIJz2wSW+AaCMOF4p8/oMeGLfLLo+Pd3Y3w
k4uNBCGGc7zubnL5lKLy/ulYFAVVjfAFRhjb1fD2aVpOZ/vOxqln1ziF7Dem1X5pOCSYsY+Hw0VJ
JSTJaJ0DObgS78+21scVWa3FgG0MPKC1WEjHtZj3ZUWQlBYxclRBdTpEU+R9N6M36CVcd8dU0zSh
q83qL3rpvywlZVo4geA4s8VfOXyrEHpsTe4vsqKu2PGpPeO4WBSioVvIvWOhU7wBguZjljqtVLmb
zJqwDppiF5fUqUDAWhlqwZiUIxmTzQ4mkZjvFJRmjsEDIdty9UNewT0AuTzRpqQbnGvahQT5vis0
+1ckGYfECl4JGNaTL7qeqeXhn4xi3xymhwPIEAOD4I8zQs6+ihjV062N8bGmPt1bYjtG5i0vEZqJ
Pi+7aKtbVKjhan2I4ESD324RoHXHB26gFy+uj51OixaNkb7s4CHPUWgUpYDrO8LjrEMJEY57Bq/M
MpF9E5FHgW4LeXSyOyc71CICfBCA4GnmElTFLIyf8bu4LCIz7kgrSOQLCvBR9uV0DNyG3wd+Qw7J
8UlbyyQ86BMYo7NjQltrg87VS+BWAxM1098xj3Q0B8UiwM24iP9TOZcLCCQLsdLTih1Xe7lB0b5U
xapQQTx5wU/wsOV93uLZdHxPIXq/1LNaxCtC86NehFCswz/WDL0lbB46YD1M1iJYo827xNtXTspM
P59PJozDmgeFC1ZSLPvF13gIkZKJCf7cp4323wlzG3x1d0cV/nvIc/73y8K0mItTzf0+jhhWZIBO
Iz5qOe6WEm3L6syRt1jXqLtuRmktIZDdZwF4x0nYBOk+Ku/DYljIcDYc8Wh+49A9InRIgqAVO6xq
+pUu9Le+TCQx5d9eNQo34kzQxlssDH6LrrNq5MuuWW9yEgEabN4L5moECCizIf1K9DFYFzNlkubj
bswCfFZatwIJTRymUMn5qjgsy5UULFEbWqcDyb5mhcIyE63enQynyYksgiKsH0bNnMhorhIbaQxD
746QIuAd4Fm9rGClhu55rHRO5ixtVBhjqoC0KsCqDP+srrz+aP4Awy1mowD5TNJH1Ebxc8zJB7GX
/bAz4zhSx8kFQBmIcsH5zOHx+G1Yky75Qzc/wZ2MTvIVwjAswb1MEJ949ADcrb+rqYIGttKk6pI3
mVXOcHxOn+F0TZIuZr8VZMZhtGXTiBmH/6YgjU9cZxe+oRTqtBom5riG7mJaeOwPXX3xctPCTNz6
wI3H3UBXpeoTzB83TLbduWGaedtonTwBfxoQ2Hp2ezvoFeCEtQIxLgEYUqRczRrL6iq5bFpIN1pb
lj15L0QD0Te64DFELib4yD+ukTFHxxfU+l7psUw7B3tYnFkMh47R5ZyjtgY7vygl/4k+onxWWey8
kH+l9iqK78n+eiUZkQUlDPmhEA4iLfHrUgpXCkvdYoVf1jU1d0np6Sc3c5zSzLuaynpy93175rN0
i1K92HKB2ObeDYCRwFALGphyEaFt1miequf2wD7HCaG0kszd3ZKJKdgaqtLan43gGcx9m7OiuFCW
XVS35c6nNaibPiBbiNJR8seMsvdmq+j76P707A/2ETb+qryUb6BqZ8VeF2WGzV+iEHrdPt9NIvVS
uwxOlGDIxhmAWHJ+aS0Ce9UG0pVWChFwXP6QhYxMdSKmfWYDGZbuMkjrDo3qi6X6VKKY0dRfGQa0
kvovDoAs+LHQJYF3htzFrv9PqSQDC4CqgYaIxUiTGGuLOska9LROUS8DwUkjmtLcuqNaRM6MJfDu
5FCAnccr+zI6ydvMn5J9pzRhg7ebZ5JyHJqUYYovyjp8ziK/K3HF9hefMTx4x3VcbvtZUY8cWN+O
IomRW+KnW6sssPviYBbbLfK5bEZLJXOI3e5hxw3Vr3JjvXX09HWzdei9H/yOhE+YZYLbzqq80Z8H
2FjVVTsNJW3+8zIKoGW1yX6aXPVXWcG8fj47Y1OUti0ASuLYTJrPM1otp7z9fQRwaCShoRB45HN5
VfLJlqIn9vVwl5sKHGghrqBSyLLBIfXN1k3j2O98m75Q30dOGdWwedwIlqsiOkH4HO/cvg3HQhH5
PR2SWp3tR+zWPn2lEDhvGN1W7DHehIsCwwgOu+yc92bA9KPMFhgC6jeZAosneeUB/Y1XmHCRbQtS
msbbsxX17/bSo+FsxSgPehYpIMWEb5zH5mHw6gZr+LZYfByuwkeH3l4wbw3Imz3PqkIJXKjZnLn1
T2x0MgBgZ1gIn72TZnJlMmfESqLusVpralXZyTJa328k4Poo1ThMimrB5SxMkQtOF7Yn911VRkiI
WolxzLAq00+6wnrClBf9l879XlsaOvE4t3B4adL7cgxnqFV5XW4pX6740+IdV7oSB3Dzaiqi0zud
IbAtGs+lDOciZjlLiLoftWq0PS+I1H6E/eH1jzebszeIRspImydSp1TNrVGjtOr4wIRcFQ5gezVN
tY3UbDgVhltP6ZJp9dzer1hM72tOCAxe/X/9CYlL0yqjmH9W+NIFU9knLWZAI8mVCDqR6C+a921S
T4+u2qQUJVDAy3/qNcJ5AsFlBapwV7bD5POzmeE1PNnvg/2FgoTqLuDbri+xprAeDH/KH0vAPbuz
ZR8m2fj8qC33FtDkLwLA6yxe3zo5/C0baKJLvqQQKfXMj6mxDyygF/7d1AYXFsIaJZbBneGxQu+Q
n49TH1W2hxqonSYW1OFM21ACRRukFmDVlfOmwWy++LYh2PdkGHCWMhNKxlvekQEbm0qLWSjLiDE7
pzQQ+XIn3MHNvu3AqhQ4KenRTKaQoGdj4zwgczZAQ7R0y07Ss+hHCoypvMmEYNXsOuH9uA59hs9O
Y0zwje4RlvqIQ1zy0v68LrGQlAGEA7RZHTeGywNykY1r4r8z1q4lunxc6zT0BitSfZpr7k3wqvuY
j1hB6OhhQ4f7+sV+v7Qc7HPU8Aef+4Drfy/G1B5S0fgMFytaeaSyrtxgzTX8d9x40fjx+Jk6HeBX
R+1O+v+CSPjwxIWyvpPGHlReXknVgBJxnUX448avE0jnAeufQb/eKPSVkWXGMtpYx8u5UQeDzbVe
4WyG0OogrFisWy/yK1ZX2WUEZGvbTbI5MnzpbTxQdARl6WyihJvWKpAgM9AXrzSzcEX4s51XURwZ
Q/eX4fpBfieDWak4HW5+UbT1ndlorg32ccRtKAR/9DKbjvkg1Lbso5o/bkSKf9GJQJWRx0eUkjQS
rrG2GJfQRNcCDJPPcDbpW/fMpn1wqasMSekPEKgDD5VUsoGdsp1XG0CpJdV+4ObYSA3OMHxDU3hR
wasN85gbCpkomEIFw8+rOFkMBiAVRsnPbvE4bDD2xWXwmKzsIU90FjfizHxkCGFSgH7fAsSOq9A5
YDKStimuKTKTPdXsmapMGM+pLHZMNzLu2HCCL92JxrTiUqI4VYc/sb6k1sB4sEMrSQVSuq0K5kAu
6DMUPWMsmdWLIufS3eb9nQU17kH/n8tfXvOcIWQNGAlBD3V3CavvWG1VNpH+s6P9dJck0r1KyZDB
k93oSLRD4tw4vnEYfRyyB6n+pTGykxpDO7sbATB4vKz75pS25YRt+tL2SLo+4OWK44mZKHjBCwxa
SC+NymgzejRLXgg6VaWyFy9DTwC3gKS3fxm3oUAaegHLQnjt6T3rCIAnMB7bIFuqS7EuQ1jsK+qt
/8FdNxH/D0e1x9y2B7PNJYzDL/7Qv006B2Q4plTmxR03qpdMBFaVgA3NzPUJOqF30Ick9+1L683X
jrcAQ55F6OI8lEFRx6WPizbz5JZzM+kOcrocc/r+hac+CH/N9LcjF6VGlCMT5XOnGUrh5et4Mz8U
0TE0CMpYIKdkm+NHKjNPXr//U0wpoP05w5jB9insw9AFNmIYJwl36AMGEYrgXuP8bPRP5oZkmECw
LqLz9fqa0SyG+LU4OL+RMm+t7EKp+R8hIaoIAh31pgj/uC522HQl9IhTenZfVMNil0ZmsYVNovji
tkLSXfvOdXxuKleEqs5R/JRAtDpx2q7XP3GTnlNddB7GfNOTlehrWIw/EMKR+OfUxytjFnwYyCLe
Hu+Du2cBkaubH/omcSxbSD1VPJFtTT42kqMNLq+PPzEVOj6iLA82uM/bxb5NTvJtZ8VDAirR4ovF
lXPH8Je44hZL+Jzd4MdGB7Dn5ILjid5vdNBLn4FnuhaH/BwH0e3CcRHiNJVL+nagmlYm8Yia47OG
ela9ckbq3lGGK8stSqTpEVmqTc4DjUDInnEBYzrKJCKnwWkx7mznZ0xremv8v+nk50NYhvIhJSAV
5kttckuJZw7TikHxHH5ZHQk5DU/WTwWiAzSXgZ98JIHqTbcvXfc24bZnvL9dB1H2D1mA656x4SMA
fdIB+SBQg3strPtjBAAEOpHR6RcUnFkfNLLvMvdCTh1txwjAKaNfs0zT8xeRC5sl7JlhWq5CEZuG
r6Fk3yfHrtuRkO9+ubt4/6q97O8I78vVrh28b/mdYbd4+IJEFkF7QzFVTLXjguXYMCUYS25qMWxT
IYC6zHw6wCpqM5uE9lB6P9VsqU1cmkM+BLjM+vfmJUhs4F2vpPYV2BoCIyBr+UUZ6FYG5SSm5CTh
TH1iwMI+y3+awFFEITIuaxj5A2pf8kVy793pBbfPXhLvow6puRDX9NzjQQ7iwKIYuUSn9oNTw/7K
6cqJbFq6LZW9SXGszFxsaRKUXfYIgH8NEBJ7qBNHCKKSY7hg6xQfDIKY+6fiQ1rwpgdn4WJBBAFc
yqp1ULlFCKuWhWDHoPav343UytiPljTlbfAN0VOjyXJu/bSrceYuV4VlkLY62S0KCyqdANHj9Lp3
7SflczPjiOGxJLssK15xVzOXpvmP2thL7i1jJsFwULk5eaU8fpKKrWPROfEBh/cBe39t0nyDS7JF
HH5LoDf3/SHsTRucKf/FXEpyuRWWI4ufQ27yE5LgMiYGb8PpWkbQbj9YeCEhfyWDUWz2dDdxb+oJ
rZyDyXckyp3puB5mtXZ7vtBBpEdwp3Jml7jBvfJfrL3EcV6u/fc4HSTUDGPnTRq15/UHU94QWn7D
lR8UHPaeC27u8zOo+gpyNu0Cs/7vFREu4ZVjLsxLDx/Dol1SQ1E2jjenNQ6zgFT/lsgT5SAc1fNk
xSF3FnVa34XatN/M1gbp45h9AR8Dyj+XRY0HL4o40BDa5EN2U3fj1H4o+IoOIABET5FoLD8VESPO
7npqKS98Pyw6SeeToh7nmKqoH6F2mtarEMcrVm4nIYgoHvnAAa0txOd3GrQuoDBcmFO55jeISR3h
UU1M9mqke52pCrvBo092iByEHd3NR0m5NR35a//nUM5JsD+ICOTKeC0Xlr6r2yNOCb20OLdLv9Gu
hRRWDApNBQPIEY7wPiP379aDg7Lz6UikRp2aulAl7/AOrNfxyxXpIv7GWzM8XXatcDX58+z/ylCZ
m1cfoXlyS5S2ID3ie7WZ6t+IPtUF5sMFmymRxE2j9vSegHnDSawTefYuqAsPtZOQXGXobYF4ZbUB
wqpJHpGni0fzxS32g/Uk+ZSyaaksddY1H3ARhzzEsULWqgLVb4C8IbrKRsh3uWJ0lEGwRKLndm5j
+iq4tUZjdjG1+I6xXWsUrO66NLSXLFKh/dV8EqU69EWPf+eKkHbLww+L9qaJlb/N6ngXVoXGpR2U
FZtQQsfE3kZOiCPooWOcJpA3XjZ5PI8UkIiH0Iusa6tpWQQS591Hyb2AUlbihXx+X0906SE0tyvZ
Hy6Z3Ny4KqmoBnM6uNpZfsxwilfuei/LTH8+bt41Bt5djnAbAs5xsrlSjXk+ZfFUJ+ZXU6QJ6N4D
UsbTTTHtivLwMpdjc98giJ6Ht/HGDl+RNkgA58UjEEu/XVBysBF6IsUG6gJieTaJvKsOQeZVBjdr
ZFF5g86at202wx9Ea1ZdVdN3EguLIVduERorwM4nSe7+hxagf4DhOnm6s7m3O1/NapVd26kA1Jye
/7tZDAMb5RW1PGHcCf1LQBvt98itbXiS+1tNe+qBxutmj+GBTf6tLhMItX3Se/jC6oIRzbwBvHWW
DEARlJ7/uLM2hlwE522lcYkMtoJdu7FunuUWDAGvUD1EJ0fQtHLTNzvtOQaBbqUdwtj43ocVv+44
k4NpXlWAlAhSQIZ0rdeyJtZycvCAGHE4yUtBLah6W2wgz5G6TCIcDznxO5CSDdQh+pgK8+Qlidj3
hDXIxT5cAr/19nxx8pXsHHUz73BA6gIVcGO5QcwFT/E37mC6vK4NFrjTUnLSUGgqSPsu+3r56iVZ
LSpArLbW+eV1mORvvjXbNw+QJaCs8Sdrg3TjmCK1ugW+hv7aULSU9Ipkht82fEON4KSPA4RKNOHu
RcbRoG5AdJx9Ze4LH8Kz0/YyUtmioQcAop59HJIW3RC4zAsjcPh9gl30YwxPpgpd0GMdL4uEhZDd
we50y6eBYdWWmUgkYA37BNQDSUxBsb+gbjkpSjkOofJKCpIrDM6LE6UXO3wU20VtYbRxdtfDrdoy
fx84mJ98SPQVnps/nWyRhDLOuQftcr4VfHi+ZGBsdFH60QCsypQSx+TkXxdKcF9sL+7kg0+P8fg5
6NShsltKObvrPRLRPz8fTJwHqawt8VyH/cS83uG6ew2hPaUOzCqvi3oSfn2EOEAeEgphgfvF7oKZ
fXuVFuaBRQMfA4CRoLR+vxNcz+dHVxsULcy8eQ5J9+vnw3puDFuXPSLvcgeyDTtp+CDgUWA082/8
8Gbkzn2NSIYPmHqizd1ZKRISPWABRR5P+JPlNA8qBz6ChKlfIPEC2P7mUjn5jTNqzsBUpZQawT25
qkO1N1tuhLC8INWQ42yyB5jguAKruHBo09ab8xWEw1s4wAHdoZBBK1Jeym1OPfor/HEPgMZTT2gc
Cw4an+rN5dtrc9ypfNONovfKpNONmHs3aWB7mX/YYYzWwNVeTdTeme3YeM04WnPzv0q89jMn4i1R
V+mDUcbPyfhqJHLtvSTDyXUdov+UZVh6qY47M0+RDy5vHJbUN0nY2fV57jYcGfeANpJ/hymWEU8S
JIEAUzUIZ8H0OIAIBjOnGkt/5nNG4bLzKEsb8G5uhWlcvoYwkiUqes/YxDyRVk0W9mQWRsBGVO8f
60OVkAs8mCnUZ5e0ghUIBCYt2dkHz37xlUvb7uj2dE+tOW/LXXNHzKO8aJYsxQpLCb0mbX5UdD6W
cocP7pnH/as5SZpAN/UdPg5B1zsoHO+bTee4bFbvWqpub3gVsXDr6uFot6ogRcSdcPH8ozhApVuD
KQFj+xeU+tnoCzynvyPWVj1xIZCOFtqL4+ROnifmgHsFAjAGI1UnSryZGEofbDFNV38hbyamAT6r
MjJIVl6rBtwWqd+HlKfpOOLmCu1WbG+OA3brAbl3aoLc40IXPm7Ost9Qr84Ja5UuG7TmpWNQpbTh
fhMGTXxwTMqsmFylk9uweEG6XuMQF09TKQtaWiL0iTlo6F/foKPs+CPhrRQ2+Xjjcc6eFSgJEmUT
BStDyWVUPWUX5LFfxtbkwxFFIIKC3Y4GU+GpjednPkdeAjqZ8Cucg00Egc43bIkExd7/KZ4n7dw4
T9UCJQXGIzeIxCsZ6cN4/YS/3Rw1n+i1mfWTodS6AIGcAyKowosq2k5np17hgWy6CJdpydcgn5Ag
HM1A7Ui6ZxL3BaophSTcLBkE/xzWeGlZ95c9hcnYYe+6fN1gLGua063NRgbtWm1tPB3HajMX0Lso
T/h5VDgqUc1Rfq+LowiVCoOlcCBa2jDnQFWV0kpIQpMVD3doOoXp5aJ8Y+nworiHRG9/042hsnQR
eFLMi0iJ/kJms5jaPJF7P20kEsUWAy0zZpZ3YQcqoZ4dlDn7Es4didI7mnZCq6DhrAoCHGEEQWGo
Wm4dKQH7KBLKld4EkZNvOtH0ZcEoslmiWTC4y1kM/XFgXXYgTZQ4GulDYs9HMlCXp1yEXy5Sc8E/
3Tf23+cOwvOrd8eJuMMhNg4NHdnJhODCt1lQtRRO48oOapi4kEgzsRT+D8FO7CKzOxhVdTsF1IEW
yZXwg0FO1R69cHbZDW0sMCknSmy0qz7GWSliP8FAWmUxmYSjFtetoP/iYU9XtKkalcwMw8HAk1c4
Pw4DGYPko4ZPeuvOTLcxkgMJUDTaxItnX77hHTUsMhCnyNsqRaPvk0h2TmmWXuylCwGMtsPS1NcA
ja2+Lt9TmoiVCrbbHrPFtkCpneiikdQrZMnc8FieKT0+/f52+tedZfKbQmfmBaGD59aUIyhQnyDv
KoQ70m/YW7EBj8ybyHJvlsWcYnmvIOG6BYqpn8Bva2pKLg55KcIl0vtV3ZhP2gfTNOb0Re9YuES+
fseTTXEEPhUiKGfc+oPJNIw90w0sIKe1VkijDoiR+ZqgrTWhpyFjScBk0/wiOUQmW7pB9b2mJKS+
0g4rU0P7knv5cgSmBMAnrqJgZEYkNQIFBw/5Vl/dhGHbP52//P0yNZvIE9vLYXsZ+9JAh8nsDd4/
cu3Sy/VUh4AKYHry9qkmhfddm+qjDlKFm7T5WbN9Pr2ewf0IHa86NEMRpC9s4bBJ5IOayfHGZU9q
h2Eokr9my5mnKPCgKjc6qorS+vVegpPGn43/toYG0KhBOnL/pbwU1iUDeuEp6zqIvDUzH5TqX5GE
yM+JjSujVBa+7T8di1NfueFsIGp0BkWF+toYizkekoxycAbU095xa/gv7ZmHEbLZWL50YoB/aQmq
DoEiE56qGLUL0vG0Jj/rHMqSmSfWhs9i+K+ARhjQewHpdXOFDhCVIEPlo/LVUaaBVNwd+kdVpD3N
DT/6BCq5Ma4VsHVUDXKUMC2LL00/vWI4PAc79sLXUYqUyj+/LtQO74MPKXV0oUjjZNCc4MYiMyPJ
BHTKgBvfPFkLtXA9onSLxvDqFhP6/D8aqTFTG+trqVpNV1P2xRDA4W/97LxUuIGIbELOG+MKiEkR
vb8nYDVZgOEbP5waaLfEt3G2/SERNmjr5XujqYdAU3lwt6f19/a+BurtRYbs2/htu6geaTEu1sb2
jkGXwfnEBNTZ91Q8SaXoSjti2l6uGgNBaPJhLI5Y8A/Uv/+tsenYvslh8yaKLsrDn8BAHSX5Q2vR
SHAkuOve2yKuqF3Gnp0Wy4OzWMVS/hYJ7R5XojLYjwdTUNwW65FE2frcwcPBT3Ldw7JHLZdpSMLK
RAKbvpTzV/rpjQe6wOG+KcL53AJ6GwKdydNsY3AQCjfGYlHlAy5pC8xjFNylWtNRvDisFJ57NuHw
59LrVTmjmPlxIBPmw/xm7y/sPkmS/D9bdhMjRQPFEauDD/ok6QShimqayArutIMyRSNDRmkFP1SP
+JbZf8zKDebk3pY3O0RWxfQllo5msZhmuNmIcCL1bXPkK+4Stm7vF7nFv8qmbY89m1CgUABbc54X
9nGfnY/eSYpDyRrEQZpSjP2ouYOKvd+vJyUoUcnlYTKR2zLh8GNPvhccXx2hKjYvifDF2quuv5J2
WZU13zBaSkLWqc/GK2mqCVd+2BR9l59Ez0GWIr9dVuRIBJjtNQ3nF9wVXzhSC7wHEiDK/slloG8j
6oKexZFssMj9gN2NwItAc/2xFalkbGnIlpsVj0B06BYi9UsuxHodQHsrzii+L/2X2L9txVtq+lKd
lAWOUu+Hy+7NozANQvj+BctBlVz4o85UFbghl+Tkak0j/BlZ6FAUcyKDCxaQx8gX4stwX/FL/rec
peLRPLFql97WG28Ky5aAzBheu3w4qrO+Nh5y1NDsGFKsKctfHsbpJ7O/1zpcsziuI//kgi3WTV/Z
ogRy2zUvCMZS2ygIeiy3JoPXkAOZtSM7eOYOvHUoc/W3KA5h3MvDespHOFSwqGzYeQBAj/j/LZT2
nGDpdF49nqqPB7iLKvDoZ0j+mxOUh/WQ3xsjdJvr3YzTa+m2SbAl2EzhsZMmrfWwnximoDMQ451g
G0XLKeBW2I0o7KMgprjjnkEdWGrADeM7eQindRoowOm7WqtlC6Oy5U0AyBvvHLVZ41tdBeYc4cwe
oHtsLZzGcwzTCGjzoyuFtmaeOInwiP9fau/tl0Zu5lWMKs+u/3IP3ARCmS3cbfohrwvbxALKlpLf
W8e2dTQBebo0lJ8qcT/NqO2oOvXITEBVQsfi5SKjCt8GlBrWJMmbIdjhw7eIXWfSXGDjV97ASj95
P97kRUippTVg4IL9XzGRJYFLNo8LZ4a47XHwhMuFbxkEQY3ClBAqNRM0lGszC7xy/tNGv0x3JnFr
6r+6qUNVJblrt351rFMN5Py3Ya95XNQyNTv1QhcxK3et/R/+w3eBWEWaR1SgaLSk3wWuCnzvEQbT
7rHDx7HHggu4NKDnmMN6U68TybW74mWyRdAiMWwMCCK8KkrhInK2NVoa0z8fx61gAUSKbMogfDGE
QjFDJcFkEcFdtJTjUYsKrSwNSfDfe3x60EzbaPB/hv6XB2AfT6gXT2sdKHUpjURt5ZGalqo5iNBW
cFOe6MdCqkO2WsYw374wU5f7B7WunvB2cePc2sUDOtWia0gF6etTo2Fo3iuH8SeFMYiWO30X+qHJ
YZ9mtiMlufhqnLNqrllX7iYTd399u/+PtylsdasqDPBlLPrefRpxCSegQHnJS1bk5xCB6CZQjB3u
VK26Lm3GaC8bau0Vmra48f9v4kPLKkPYPoSZoFMVSGalCc3d/gCYFv0Rf1rTh1C6pBWsiEtBOy28
KyF93GU0fZ8N6TO6VtPk+t5v1e3tOePcAJJDTXDI6FvC5X8wMdrWdxsvrWF8lyhuJ3IaOIITyzzZ
qNTmTWu67GfP+7NL5u/8aO8hEJ4bca5rp0mUwqyYImeRYlYkAzUbGM2fPEKJzSNer6gQUUrqvMjs
o9pK1ThC3b8D/1Lt2lK4XG2kvfyWlhHrh1lVKsixhs7T53m04avmg0Lc/h0Eglp+fkC23ArKIrRF
lGM3WinI+fVm7lUnijqR6vmoY72Uk9vZtytZxKYq2togptWKj1vczibAOatwb7wjR/ngcQNchkTt
2/WsgxN2YnGU+40Uu0vMpCMVBbdPVDqI51t2bfa9S8bvJv7Dc4FBl65FWpATphwBC8f9/Zgd4Nhi
EtBHbgCdG12ZwqeX131jR4rcrmd3IVwqsKDf3PIGzF7ONVXBXcp/6GVgEQF8asTaK3t6CfdluE5f
vOi/9nH8gbyVN6fcBx5t4U1DXF5NRcD96KQrS6vNk8HMEaUt+xfial63o2I0LkL+Y3EcEGd/myzj
x4Ha2y+O65MXkf7ZL/uu3AYs22XTxRw2TANDzlTjtOJkfnkcuOBZRvcxYArJJL3eKyQi8Jrr6px+
xylEfoV9n9+SoWlSQYHkIe++MwNa1k9gAIC8w9/2nebLn1kRvkbk0SUClSH7c0rlvm0K9CEwjzaX
IBPq8i7Mw6E3WA8Fta0/v2pg/W7hbDevNlpFCqtpL9zrgn80Z6lBhJ817ARlfkJEn+71B1I0vJE7
eXTn/Zoevu8Fe5vxzMEFDWjVs5HmPoKy7J8oKZvwQns7iqjoQmQ8uYH3725+t97R1i3zVSaG6PLH
ItFK5kMzXMR91x8ELp8V6KyANRXBeJDDz6D7FxFYb9esohkONNczXbOVw1venGlD0z0gLGeUmJ+7
8Wz6Tp3o0kYPMm0AYUG+YzEKLwNbhbtis2M5TPmm8qq7f66KCxEnkL0EgPSYqoTbPRv3ngm8If1P
d4/P8jBICKpcH6w8qfXNLxscf1l8cosiklhBtaijvzwnt3/8Xrn2pw/maFQl8nSKb3cNfoOlVUw3
J99u4/LGjIvPJ3WULZoKspZpWZUie9NE8MDUxtFoWmdBTMBQGBz1DPHA6DiKLeLxQhSlNRB5s7T9
dcO82v/q/k0aT9e/ppbNWIhl9K4PWRzudiz5hask92fXEMmDT0hl/hkn8N6PsxSLhQ8yesnaJ59o
NHZHvbyiEKhA8fQuF9AtqVtbBooQKEMkw+IMf5wx0jFhD+y9RUDVWB8wVJIokotPHPJYUS/sOsD8
Yx2G0FJF+Yl5iXRfiXFmZqhap028sK7vq7apRSK1rZ9tKm8QaZGj7oDm0Ys/QP5HNz77EvXKWvfp
QW1odmC/aCIGWrAMEuSncoCGMGefmh30AaW/544BMNXlH4R7LhiL/JPsgvtT4/SbRIBWdNaUtPk/
owBCyms3PkPuMsH6yitp64Te1aONbiGtvTfHRrv/k5g8s8rfvXYZlamH4pZGG1xcAewXJcOW11k1
4g5ilAVjgQMcT3z0emWAYbIiOrCH829TAK99gDrbdr29F7wlmgO4Gp8J7DdEKaajzyna+HIku1AG
Rvgn0z4xCVX3huu1No2S7O50cehteZ4UErtfZG7xA++I9jikdlcewCMuTcZAZPPmHLg9u02R0eP5
sr/cidEN38ZACIpA04PwFDQr4Yf48ku/EU983A93uf3ekSvaF5wtKs8pRr7yhT6w6B2KTd3BMoMH
rJALE5u3SJwEFswtG/0AvQRGc5mJklIqD2jpXNs9VtUTXVIow17QF8mG2bxjgexur8Cz4Vqmw61p
wdBF7FZ3SBndWbSxCCCDH7HH/hnj3An7G4jMdlcIVDmaHAKi+1Au8wdeI8Ce/oBzdyWQbQq86h7T
TxOKBea3eZUEwOg5Lj30/hIpb87BKl+qOJhJcVF2xM7/luVyih3zEcRUS76QToq2Oq3Lv6+jZDCN
T+OEWT1zl9KNg2zg+9wMS+DuSAU36MFVWxaFGeay2cxBnKxhp7XSsi/+usLt+r5cfr4CCMqu1Y7j
51fpdZ4JeU8fY5cTrjcvDKfVt2m/Ecpu++hgXJ6IYDNIvpVk1QQKcPMqP2sSQ0Vb73QxoCWqP03W
jjy53IlEshCahZieuSc42qOrMXgtW9w9eQSHLEcbjlpvfGBhh/w4t5VMieKJoRCnIZAykLK+46HZ
QORIfpVQTAaDr+WcCOqLajAI6IiRqIFVBEMZ52VQ0W4725+1HYOMsXeVvwgs4/vIv54fYZWFIg3t
xUZWkY5TeJAhxAFMbw76D6AKb7Od65W0zBsuQp2vCw0byaMKNttjo9ze8LY6miDgrB5dKX9WuwH6
oqvf5118m4Iefg7dGx3ha1k3+lXK5CU2AogyLWvD3789KwaZF3IKw5dBMxJYHuCe1jOIFJUMOXFU
5J2mvYwS0fAB3CeJtYMz0VmvSyLlhZlmhygyhR9UMuHvwmZPSd5m7mGcsrXMtxmdQoFsFsHX5phC
U+gyx2Ax0Xrt5t/2/e2zCCttWbsMXwr/t6NkyYJvxyfH6Gr2kFrAkcPu1AP6Jmu0EMn6MXhkBjHx
0ZsBh6FJTY055Di7YWt7V6r6aMO59y9XQq9QlGurJgrJ6TmxRAyt6c4BStSxJWQsN/PMc3lzsx/f
vq3n6hWaHOiP3p/k2DfrxRiJKts7S0xtybpicHCOszriH6I9srTvkScjaVgAfsEllQVOaQwM6DqL
WkYN32exn5mlHxmOUZYHrOCY5q07yxFDKCis9RkD0CvC0Ic9YFH3OlCSDHSahNwxg+L0q1DOssH4
b/QyidqNpBzpe754LIix8QyR+6/fGjyufHIh5Q0EulXZb5smt6FOFyoT2/hCeRW4L9tdU9G3Ig/5
GQmy667KbKmZ+vK0r/gkRMp3YfShGo/ku58xQNovSYMNEBXIPD4J0ZEIlAvxi4d5KlO0MFhFI5Mn
9hc0fth9sId3nZEAfxT8b7S192MIyigujI10QQNLqc0JphMcFey36hOxQxmRE3u1nfh4qmqDjmgN
Uq/Asjran7Rxi4+3LniiPjZBp5B/5RcHAd8vrdQkFjTHfxv/Z8H8fVW7JIJAjxgj0NLlLgGrpfF7
Esn2jA77Bxsb1hus5Ho8GmtPsL3TZeynxJG4gqvVHSaJkta4UkHiPxnRG+conrTAd6yh4PZ+Gd1C
X0AHE3P/8MQdZA/JlTQ/q1q28AlSakiHoIrAdi+2ezEWkMKez+tyU0F/r7XhCjkGf2ucT4a+lkER
9y8QGDg5f03sCDNanUdBytV09TpM4jYnsf1FV5NotlUTVvQgcAFr+oN6aU5kNl8rtSxZuuG9rlPg
F4SIqpLFhk8lT1/ljHmqNGrCwo0A2XgNOntlck1l5vK2zC0jJ+ZZRy8MTtTSKr6iOpOSYwAipUQ/
de98Vd0i/1U8L5SAVHswTFgVlG+/IFc4mSE0X3nxHaWisIYSmbkwkRK1j/rabP+uefby6e8FZvp0
Daf+Gyy0tUNE6P68FCsVrrYLwDfKF0OAzHzSmOddNYDM5CsB3BwEmmfvEYuxRglPG7al8kq9jSxx
ybi6AERcqZVI1knKlYkQ+Z2B29np28HoYdfoKG4+SLHTYR2yNzPdi1kdJ06mKNeMnRe69zSBftqm
UFG3OZd68T0z84HMiCx2Bndz3F+KiAok9Ma3WHKyEERSWN4lFwYKK30N3HEGKu9lyuk0/GGInnje
MWDTle+qiUPDxAtmKsnqUbfOBBK6Wr1fwVTSDmKRXrq9xcc6ey89LY9wuanNkU+gHzy7lrlE1jY4
bgTvHs62GDExtQRf5IZ4TrhdKV8E3IlKOnw6b1T9rUYYGoMf7nKiwlIwtly1j7Y21oxgegTSsCMt
WU/D9OLgvNMpxPc4lv3Ot0sXI7J4m6LNz2zG5xZuGBvh2+uD0U0tHR5XwlS6nqpNIc/+lx8owAfy
TzTrw3vMY3TGb9z8i3QWOFDmViKjSuN9qa4hp9VHCusDZr9w4Xs+7gx56iGdJhGHtGOEuzxxP4TU
lhWeIoTWxcurEfjTkhVCPJlMaJ19dfcOo328EqM9yvIAj4Lpx0ODpQYlOvda3lUUsTbQaeylwNwL
ENm+aFLOnGlEKqKj2ne7Zu3K2b33wmD80qf9u6iuzxYNGO+4AR5qFkeLTEAjZea+OEiBrXjY5Oa3
1mqQ1iZs6SGV4ko1dLVtyi+5eHuIRqGYWRjudiqNEphXAMV6YHzuxNUChyTNSKVg6/G5/MS+O3kR
ohWBUGSEHmIPwTFSXWo5x5fzLVDN6JsKuVPCpdIAQG4SkK2ke6RbpIuiKmIo9XOGkiIcAueUqcPC
1/KCEZ/JkOerHlrxmnoGsYta0V5wQiTH14GbZAfQe5VGiOWx4Iic3swlYJ00od8mQfYqDaAFhEDW
GO6cP87d6ZOjgtHHX8kugbUPacZ65VBNQV7uU9Kse+F/EiC2ncCoKhTyRxce+n6OLx7yTmVvwX5L
1CMr05uaRY4zgE2UP55pYnYFtJLTRcGsxPKG5zRY5fzFGm+6kN/ZAJP5Zzz/oJev/ZikSw4ixMMG
Eh8zSSYL5bouka5gGGkhjDp8PWQRkhvaCj0/9Gp8dFQ2Vmv2jPi4TRYOdCYebAMe8fWPBfR3zdN4
zAvEP3icgewYu12bX9QyGrz5/EvtjDQOfLGedWJCq5OBzLWU0ZIgJ0sWIqu/eE6CvnjgIIvvEmpB
sKNtnOR5HF8stl3D85As/iPz+w3Qv+KDZtxevEAR5WbFuDytkIuR5uijg3Og5ICupO8KUm+JLJv4
qogUcbzBTTXHkXFqV91PwQCXDaK4aQTmBGx8o8Fw5y61dLFJ92g575IdzDM0oEXCNm/YmYAiXSdE
3VxRJJrVs7vpOoxkJakcexVVoakFVLfZpoljC358qSSkSmc7fSKJmVdPvMxBIPR2a1dYyYkzr8qU
QBDEQ3PXXn1hBiC1Jxlrk7qFY/95TuP8GPgp6+trne3+4EfeKOOziz5OvcI8k88+dNnfsX3mLfkE
hfOyuxefz7o5XcwdSJ2uQo2RYtUGJyppz/sseLUTVmycaQeZ5DyR65VrPpkRJhfnECEOe4iLQg34
6R54Ew43q5eB6WoBbys1i6U+Mmg9hV7F6KYznx80fht2HvBTbRYZZZjegrJ2hPMi5oKZSO5fZ9KA
LOYM2SKHRtybp4yuiEEbln20iLUMmgwmgBkMKmw5pHF9j/gxNza3yDH45AdiGdJcd1QNfTvWW72P
f/2nIcQibtd7P6ynC1J+rCFwbXEU6vgvZV3Y9JJ7hdkKWZPZP52Ba+wu7EPWm6dyQh5ZHOhjl89F
HzB84Q1TcTNOP6tZGsXzNBNv6uE1OXdJsPRd7guennh3O5FTTm1UjJrYCDA3cOyWyXS1k/rp0iUW
D1xJCsoWjR92pRnNxjCGomHhMC1QXCZxq0R0tGO41zMtiKiku7oOn6Xn/sncwn7ntWmoIQfOd238
Un/nZOQlc9G+05WGN5KGO6uzVtYUEIEtqCBj2ruSry8EpApedRtxo6h0//CwN7ckQxgnoLY9MrP5
NyQJ4WF6y3wmUOxrP1n/RNrbLMKQIo/U30MAh9Y0r6iQoFiYYl2BQpOJioEyKBIS/xgXK9/uqEaJ
zyBNO6lXW4dCAE/9w6QgHfpqM54JDzlDa7+2+hu2zkJOZ6CVP1RlfzKIYTfgRIxmyiXf8zp6t92K
THfZn2vF1JzMOWXeEMu3KtDT3pBAXoBq+9+xGHZiw048hYxi09ab4qUFiF8VWyn0pL1kGjXTkOHe
mGJQAg7ZqZ+vU6AHnvdE4f8RAbjMBq6foOCkhGPqFNQ+rxUDmmeH3ubb5XXaIOIv4nqsB9b0kDJy
SOs5gZ0eOtCL07ewagMIsF2OZd85cLQRhMWbZdtSmefO8LoPOg6rxJhvPr2YwYLkmqLHP0iI2pqJ
MTg3rl/Sh+FBspHSvzXDpVV5QtlN6wgnSS4d7K3ib/fHWikh/MH1hqxMIruhPja8g5FLIxHhK1N6
iiCBEVPp+EGz5LRZ0Exq+iWJpejtQx3ThUEnVtNRGX1J3GhdoklHEMMwLp+ySXhcJK57xaggpl+5
eMVUWhIqZ+rYORKJJyTc+MHMvjycQVJTIB+8SD4+9GzT9Ht+NzMHP3Q/iEr1qaspLScdAfIB56iq
T4hcLYPW3731w90lHRC2/gFauVDmQSLvwVuWVnzhmO+aVI8MSKSsJluEbrnwaGoTR73cn/FHaDmi
QrvSEmRI/EZ1uX7+SwD+hnSg+yKeJ1JWIOuoSMf7Ce2mCskS/0cenvIWtbOg6H4pr1S8mSH8AHhR
jpVcBFZPBlBmX5MQLTivfWoI8zdu0qSieT+0zQ4r8PxWfUqn/I4YTrGWD170K5UsNoK2DiwNLuU+
EaGwv9cnA/RAl7OFhLgvPubCY7qm9G8jv4jXoeg/RcVtLvDUmeCtk2trRhRgLYnWgSU078dRuzCm
31jrlXhvQIoRV5wuZv4k4riYKIO3uE/5oFPd0v7BS/JmzmcwohrYo5scmMRlvv29f+ENHkamViLS
XbCi74JoxhdMUo2GcLgGWozKTRAuU/Vo79UPeyQU/87NnDpf+037Y+gv8GbMMIAq7DeZK+tegOZn
X/ZgUYDUT2AQBuVW/GaoLAKAdBphNCohVTh3nWl2w80cXX+HVGij5XT4d3cKmNE0wpp9SAIgixBJ
YUK7Pdkp4XMz2qofqsF+mAAEZP6M6hxNMqIPhDJZVf+jg4RoBTQ6PYqnK2/ZEMdbDEpJz/QCbrwW
EEOq6VcakihfjF58qIhZJVBCgkj/E568fAWZusIg5GvDKWREJL34PXqZFgApnWNMU/S1638EgEN5
LiX8cC3+JlfKNDEAnfdbeHYSH+52nsGKEcGaAsTj45wGUAqm7/x3PDB8a3KV1TbY4r3O/wj2LCGK
lgj85s2dGGXRe+oNybwpYdNy39h3qpnFFPdPQRzhkZLGbifTD42Q3T8SJbG3MJ49gg4eXHc69Bat
rZPqFzMOMifOHuYuhdNTY3MU2QnDdTrQx7XAL4RwvPxhFGCdjcPDNb04YUntCnVb7OouBNh/4K71
jpZ9+KEDyeHlLG1b76N6aY6FvS5737mWL/Ls6a3RKS1utx74VLXdzsbcL2o0jdjWz6VavdbxstWK
LEiPnQ1wTe5h6NdGm0QhBJ2DmwKK+E6hcpx9e60cm/Khrq1r49zdlDkvRmPAojZeUnARr4QV1b5P
ALOafNPfpAdwz8KYjjzgkkcfYmNwW30II+gC8MxfPL3A8lQLyWU1EUcqLrhA8aoV5g8GZas2qy7k
exmceLJS9zFsPhy2ySiXYgG7yQSLR6VCOAf6onrxQEmv9zeZuektxf1905PH02NoZ5G4JIA/vbWP
4wf53KyAXfd8dTa0PvR6axo99ceTdPxRvEQcW3LJkUtdlI7oZF9zRbZ1DPWHspll84O/EwtjWBPa
6opRRIw395IdTzAeoQW1x+U3XJH6SwMMrBmJUXjkkZtXnGE6q/vS8AlbKOpg80osNTicZFiJpAHO
ba57DDu443ilyPzUkwBBcnpsbNg8VFW8SqaV6tCMXMqijDIh/+Qiz0492DCS6dVR1FtFbVgiTzpo
0SRLeSsXtDHF6eUU2VQPaFhDHpin4xZebF5cMAPVOr4CxrTxDSFaTdCcnAq3+8WFXHlsgJNLf4Ey
jeC2wb/QkWslKUVAmz3+7OWiQ0ZdKarF7woXon4b1mhxWDgYxdTy0RZ/GK1tnXcr/mnbONBtg/fi
o4a1io5OM8P9Eh+9Lfuuf4QHB/C84kgPx0Fd4C48OkalIBllEGfNoFwvuc0u4fRuDeFJgkVrt1qU
ctHTgtN7DywNdZPNuaJ44R+zQ+UZehpwkuAQCEEXOKfCY7+g3Hokv4RSTPNGTOmNBrFC817P1T0f
OncNAsxlPyJxt+cPvkL6G1nZbBqFpJoz86XJOZy8yA7OU73OQvxKbmBuXe7vaxO+WUl2y00oVoCi
pPxnu62JtwF5fgDRx16Z1QvTjti+W9ldbLF0gtlccN277eCOvpkEcoG+ApnpaKyHawN2qgmic6Ss
D61+D9F4ca5q0Z+H8hHHGv8/bGRM8CUoKYoPC+WW6MNhuObqBN2dBOwNXDZAR5a2NLereAUV6Nbp
GZIGZggzvp4rOhx9p7IX7yEOAOndXoVqXB/6jq9O1yJcz4QIq82EFgmW01o8nz+GVlcot7BlaQDO
T1MbalZPXGZxRTrRrUofyPYlVpTe4kf5sseUclLZ2vMY0WKOHcDSgncb+j7POKy2MKVVpKupknUX
FpLHovCn/VJvhVt+9rYa16hZWnDgy6aCBLM5Njsrq8s4muo51SQAfpTF0+4zYFEBuu4cFeQS3Agy
CmDOOwWTHRWAOU4tJHnJnNk9HSx8G8vyeeNzBFXtWYLOwZLzvIruByrgK1HIRh0cp0VwQxDrIsv0
5vlHZizGpsFeaZSaYScAOYllxxltpUrYVcK4p7N513kO/Ygz6YhYZdk8gy53R8ehuWKenOzGndjn
4GmoXQ0ONjkWvU1DlgpjFGJ2CCK6DRtNPtQS77l80HXowPUbllzCzQyyIWKJ+7nW8Gl2pxelYNxz
wiIKApvAtqU8OBHsxbW6ewytYTwWD8A8TQu82Ge4xGGM87xWchqt1VmbF+tMWLffXsJA5K6ngl64
mCDCjEWSuDGlUx9qOwCxInnaiypb+eroZ6Y8ycuHac1ySaHKFrytxGSeqFGbWTrFnzDb4N9/T1CF
Dst62taEB9QN7V60zEuXDnWoD6n0yoM/YS8YN1GH3VmAPHNuShW288heLtaL111t2m/orAQSBsTD
7DQ8bWe9IPOmTC70eok7p93fRh7wQffYPIb0SNLeGS6FTHgfKHamd1zmOuxX7pPYC/S/8PCAIJmi
8Z9Uk1rgzYzAlSV/THqXouR0btJioNEDsBlMMDHn1duo3bofdEvrIsDlmYmCYF6ZA04eCZ+rWM5o
s8/c9AMKS6RZNr+0FU/wXbjz0osG2vbzbgjoZwdPgxpUow80CXbb9x6jCCXr+iYA/jb/q9ldgW4E
Mgwqkifkw/ZW9AWGoW2QZ2Vh8u/fGbJq9uwNEbZ7BZ1o7T8JR0zBe2DYP7MpjcsSTDXouke7E5cu
TjcZ//hK6noyiUNUum2dnFUja141HFWeNvKbbROhE6PgcBdZ5zf+1q01NYOC3UCxkJ9PvvtoFsKh
TGw3sxxSVrEhKPGnMBNvuI4CzMO0K7phyHkvLIt9LFf+F9P5ufOw4uh+KZF+RgixARm9gbD6VYuX
Z8ocKvl3QR8JiDNNCX/62EvKzRMF6OSiXDAT/4c7GnCz4IRF8lrtezZDZKZ0Xh5RqU15Hzrt9laA
R5FVv9qbVtMZDgUqcSowso0E9xqFy0VDPqfzoVtcH5DcF0BiNeRVR2s6hbhSXhKzJLyHp9hlZPZs
U1RM1SPOll3sDU6Kbz/naCxGCHb1QH5VN+f07ViV0dMnpygeyxiAnY8sT8qF6s48RitvoAHkv6Vx
0xyp1az00rpR/UeuNxuKxYB5S656d5xU0HFNnr8kr24JNtgZE3t4rfh7j63nofCIHWIDcn2salpo
Q4Kl9+3cwNPooPmD2nknSWBtZ4lBZGxLCs5v/7Ic/wWBT5Qc+Lns2s1gPG7EHBRyJmiASws/f4+d
nK9GQETq9/Hk3HDT0ltSM6v0ukUIiin6veFgkDpFkKsHK6NeTumDrrIt2VBWxfW/q8r5g/ujZWqX
PoKgOEFgm3ZeX/nSQFNoBFFvGSy2XLXegQeKskcuxV0NOuOWTGYAj3Nz4DSB/p7iCCn+E6gui8XD
z/2P02XmVFc9EoBhAZ2RrrTqF3y6WrMV2lQHe50W6+XrILBtKqs33T4Qd3IFu1JPzJnjPS1vG+uQ
qaXTUQlVcf+Brn94cifzfigVKUovSUReuIWxKLAmRrcY98KCufCZ2PC/Y2+VTGwcmtwyoD2eD1NU
1XP8QCfZJBHzBR5slUhtuIzsg0KSu//3DdywTn5zyt+HwG/uvpsWTP3efSEAEUVMs2qc8Ejue6DS
B74z3sqANQP+PLmokOJw4+BQIWLfY8RbtseFa1fVZkITMih3YKXd/Zk+NsxIrigxgG8yuxKdUU5V
MU5svoTn1UtuHuJQMh5K1DB7z4XyRsl6Ma+zBt0EDtScUFkOEORy8AcROCysZ7HCpj41Z2H4Fhk5
14JeBUzRaEMpsgfIPh18F1qlExrOMzPJJmj4c6qwjNmEiST8alW89K6tte+6agdNAAr8craGqQ8x
YMMUSox8vXJOYZ/jLyg4ADBTWlH26vfxch+BDFkfPWvkOSq69uIvZhxULoOA53VAD1qsVWijz5Xk
HAh3XVd8buDIaLfc0pkp5e5bfx/1U4WudtrzLLJ/KDwKjdTu4O/+VXGrzm+TW7YnwA0qbONa7NNN
B7f8V2oBvU4Qg3Z0uD1MXqj/bHTqw6mJWGSPsI3oStCSXJYl+j3zGvS+xncmi28+EnhUAvLu5vtE
H49i/XEiay+BS06hmgLTOfSwzUZnQsZHQ0z2Po1pdlkmtlP2gMVr/lxmMHAKvz66luyFEQV/5SFX
bBLeGPVznIKnbUva09sKxptfjFNqB9Tpw1U0ki18llaB1w7kDMoFptzvMozFmY5PDa34k2m3dGZh
L6+x2wEJK8qqGx30FuerIjnF3M4oIOWbTjzE6uD3CKFMI8IuUC009aGB50JCQqm7haMFndjSiA7e
0ofQH/3+YQpsOrdMC2EGPx3gJWMMs7PhnKeM0cCXsrp03vWRdKGJfxo9FJxvhyKaOO+Bs38wCk90
1Yu1kCbDdLparBq6rf6SDvB109WltMUZ0uWCMwY9rMD+tol9I7W/S7PBL140rtW/a+MS/Kv8Wxf9
l5BimUpGJQbZBWtxedLnHBTYdexlKyp0phayWPX5yZ/hBaUbc1rr2CdH3fcTdDzByJ2uA9pFi5A/
1X/HtOareVfmrxOCWwhAZK0hu15d3L/O60+LeXGEeyxMPyPvNlCq8qIT8078ck2B/1zqzWEXSr/m
ZSWdrJs2KUzQwewEPlJVs50d1iPuCfj6+xs16xIPyepIpzjQedVIW5YDTR9riOzHKpJgge2O3BCl
NtYjvHT5JIp7m8UyWVg+kYtUK80VRGFTFxQPeaf4ZAKsiwgNOitpPeOApuDCzlhtjAX+rhOVCRZ2
1trEUlGYwBSBM2B12MHDNnpxf7MD/mjy4x+14gw6lSIwk66KcDwQ1x8Mub7ELTD0cQtqDCXUigfj
J5se/DBdGIW74ycs5sP0EGndsxpePyLWtvKKzDDH+6NYpNzs7GEt0/w5CyCxG1e92rALfGeMbjAs
njwqlk+3RmI94eMYAA3fh/+ocXDC7mPh9JxJvi9+QqnUEvtUr8xAGwrwlNpXohGaR41gdJ996VF0
QrJFg3qJavNcZoyr81C6KdBpY9DYSoxmXFsuwNBY5HTJTZAbJO2bmK+OmVXuy94tD4+6KBqWZTXJ
ar2f3RoKbxEUcnHESl9OK0fg0xBmVnPnJLA2uP0LTiyyDJuQM7UV/3fBsvD4JAnkFuvANeo3FCBX
2YCyD/mSUXUNCxughd+45wt9VXoB13JFlRzOND9+qBjePcpCCOOGb6mxu4JHOs3onrLe2QVtP6Lh
b8IUuvTwFqPgBd4zrdaogEyJfeQoER0jbQ3zTqVsiZIVQSBVKXvm3DL62JzTLnxuTXsb8otB17RR
7KFJ/ivQ7HSItynXBHmzY8wjH6umKy4D/zU2QAK03WB+8L7lPuJEw80JblRpZfqYJrA6Kg+hOsrR
jkcThbSCQXT517sBfpiwrZM2v2OUHxFzGUf7bJuMn0RUXmT+nI+HIqsW4nslHhrHu22sXITg1qqD
633x9yYBd4Zmg1iK9PMlAOzicPIFnFizRRXJDP1D5TdQL7W6kF+/l4FTWhDC9GfdwlQJHtnQZsmB
tJ5tgf5+7/8QuM7CJfc/XDx6LVU0CKeOZjSlnI4R3RfTAM7uIQObQ4zUWyQCX3es8A1cLv890FLX
6WdoXyiCzMCr9zKKzzVcJx8q1JMltk2pH0zIad9kBD0c77sQRSAUO3GY6ycgwnZZulXyd+HV4fPc
R5oR36nfRsAgGSEWPXhHa2iBc8Kq7YF2lSGqQ/bi5LUBeIfk/u2zWfuCIA4gey5RTZDxg6e/ieQK
IrjAzGgQ+ldwipphrGB51NbVdgMo5eENrkaJ3fMCdMNAiSTMx/4B1mASs3ZrBcLZaRaMnkzxfVS6
eRlN1Zxt4UoFu4yFtFQUQ0B1XAjbTScSEiBSbomt8h9ezgFKD0kaPmJiDUstgKFw4HDuOossvXk9
ZiQhgjJGzWkws/jP1yWQnwQrUM1FOfKId7GwZadioZGj9RBqqJcXzFW4dDB6dQ59RT+L+5pgz4ig
nQNJv7brm8gcn/WVk25iyQAXR7lf0UJgzwQTEKO3FgPEcRjSHAEA4RYNN+xeuz5Hxma+aG5cYdBa
ofvXnvyV7ARjqQuo05Vph+yL7B1wn2WDo8KiccOND7sb3TXAc+GGETTW3BzAK4qLlfK/gfaXsweP
fC8CO76HPQvwludclvBrRmWGBzBn4EaJDLlFJvrnWiznBcJML7nY224+hQT9IwRlvIQE9rzNcjpd
BAbc6DZxnujWyiLSPeX24DJDRosnNUtugtzcFUMp7jK5GsZ9fS/ylU/1iAm0hvUYYOg+Ok27PQnw
JUm4QORGDMxAPLPvdvVcmJpzYQ872x2RFjh5FoHdzzanmC66tQDmVf22phP8AMVKqqxi/k3Upwu2
QBPbL/3wXVOqJK2kwVlPlJ2AHfheFxzhDEJF0M2aGRMX1LtWevsk95G+HJSesQR/DSpDm/R6IDbk
/qVw7do+ZKhKBq52NWhtVOkr/QW/dsKuWnFKhWxfEyGbVfjpBWRkP0qiK72UrrbAcSFJctyv79fk
/BMTMs/uGOMqH4HrcqFTho/wPbameJol9lFNexT2QoVeum1PoAJOaoUdwL9YFdYaUDCXqKLTdSBW
/MvxswA6hSsVkwDac2SufF6KmGG4h+6Bzpb4rOR5XsUoCFe7PYxZ8a+Tta/2WWEd22xoGDncVU06
7Z/uvR1fFaC5TL7kGqCxQnS6lo+CDDBekKITEYBPkqy+tGUfPZBC6TlBCmPpUwc9rNOT2IsXUcC9
5RtH9ztIXKg8cFJrROw/XefkSFhJjYQhzWqesquhq0t/cIhJFtiLX6KGYjA8zHQ1Yn3NTAyZezbm
L0/lbmsqjgL9UKKbi+N+CITkx4oAX3doigaZflfhyTxNHDmFPJZfrrNtXQygj35vMSrPfLSEi6Db
7CK1PguoGpZ0WqTu7e3hQKVVT4Wpj8tYaCwC4Six6CTRUTbt/OV4cDbIndeJ/RDHna5XmiEhx53X
aa2NkTWwMkQx8WO3Pp5G5ls5ey3xe0UYaGeGzcxgpb8JMg5Ljn1JqRk1oUHtP9Px143PpTG2m9IG
o3we0KBZ/tg56p+/HnBsJR00Ax1vATlczC5nNbzBU3HpSklvAPXixLJiGCDpAqRI/O77paEcrd3l
43vi8mskcR0KLUPrZXs1VdVzv2dOSl08o5T1xDZIeKXOanspmnIllH0dty8Jb0spW24YdV6WkRHE
aYh2LfLwnvpfP+kFFw+Jiq8FnOp1G2G7p2lAl9gQVYm/8vWoNeqRTpKsdfSkVlfuBZ3NxtsrsqNm
PExnZZiCV5CmiKnCu33OwV+eVDEyvsXHKZZBVaQ7Nb1TaZ7viKVDHqo948PfoIRgIYwEOdD8KXb7
t6taVxRU/j4bdc/bfTT6O4L1n8bT83qgxWzeAZyKYixhPYTYNdkHw5BaB4cFuanfqEq2zjF2B+TD
YxYFKFzOJX4DufVgnHk4DF8j/s+nEB9eaXLz+kd9dtVVI9DnAfNYi/Gim88vV7Fp76BICXRGe1vy
jYtmKcmb40fDLx04drPFVQg2TU3rsjqBoJn18463wAKZPhc8r6DEosNLq2sKsYL1TwKqBDfeWnCm
gwi7nJTiyNlcvisQmOIGyfN/7peWMKrHkS3qZF3s+f58IvoTsjhNgj5ESrVQ2foBh1wjulvdQHZ6
q8+3yBej+iav2wSULKyuJ/4i+v98LVDJ45fBH96zWZGm3RtCKEZ6O0U9P6UgwlYnaEIJrlDAB+JQ
T0GFLxgttkpm5sxtd4zfxFZH6YSzdhbdZ9QEZS2XP8ypYESXQBA1utGtokTMOEnzBQC8lbGUxZ09
RxjCRBViOHY7ik6ALvsdcjca8T1g0mKrg9e79V8rn5g8XkR8/vXGtfr0Ny1gX+n8NtN2d6eT2mB7
v8QQPWGpWRXjELnJFiGOd2dG/a8whHr7EgjaOuImKOGU59ggDH+apzY8gPWF/kONyHzdE6eVkrWr
lYQnlHF8Ckw07++CjnH29LSeE7R2UoBXo+G2Slh2Ct6C1SaoXZWC+yUdOdfZbLS0ToJJYlujRsI3
bEpXozD4J//Z7fegMXE2JFqb0fQfD7KznZnxfF9GISyhLLT5exlvsLHF4Px97qgt28CWQ7NdQDXP
7dGjp+sSYuHKgBoKairJd/s08YyJbAB107g0A6Qgpp+aZr2IJWKaj7oD7jjGLnNLCqLi+/ZiZbeO
BcRvJQwWYzCafMnh27xJdunosGRx3zTYoA4KFAaEV9NWutaN6N2NpR5tBEbGAYA/3Wm+CKoarZW/
t4TKcc9sedGqL6V78MhJPsY0HISz7W12Ikk1kYFJvTkqNGTfGNJVcDuxSDBFLQ1idncBk+wlEqNI
7VB0np83fuH/GTWMICt4qtXtw5imgpd28y/hHsmCW+C42C9aGpcjHqkjDUySMuK/GRvi4SznynkK
StyirmJZwHADkinbyHsYVKdn+rFwZdIJh04h0aGHMZ8IWWbC4h6pDqUuzZfEGy0MLTp+Mm4Sr+wF
3r/Ry/eqOQKKi63D9L5A81Dp5ugNDLea/12gvSa/mw3x+hf6fna1P/JuS3vhFvNiXtaU6QKvX8iZ
6tLdBLDjFjg8fxcuh0yHkfcNlobzC07XeF6yGe/zQLdAVKI5POSOHUmQluh42m8h74sLkKT73Hia
wBEjh7bYkcsgKt0D+Y3NadRL3MtAHuWzTWoT1f5x24IgBjXe2F53gAiUUnOIihtwyeL9e01Admtt
8/IKKmoAga0ZpmuSGWYj2MhMI8ErKriJ0+vKWKOau6jjpjCjWfT3tzDRIZkpNDCRXOupYtHeB/7y
57N2JE4ZHzulTom9echqPhPjSfsKQF9no5NgcsnbYO/uYkF3Zne33620sGttq+5r3rOOZTJGRE/9
EKaMs+q7PCJYxcIBPKCN38ED6xNx0xFKDf6Hyuhpq+hJazNP1h33W6XtdHuElstkeIr5bV2N5W3U
ajlKMDtwR5SViEgEuKB+ySDJViDPlYWz94W6m7+3poFK65mkyCNn5WPPZ7pDk4dfoRKXzJpFN3HF
lzDzKgU+qBsVQqu9oiDifhFA8/NEmAjxMkE93ruoTLhSeQM0J28g7B9FaQxayMkhLccqqRhDL/VX
9vmGoxS81DZTWMLDxOXYEZPv3c/beLGHgMUTlHsNX54svIjYuK/nPPvJgWvrVQU8WfAQcO8VA/dZ
G7qBTg7P49+qJJy5jMBdnAqYo2K7WB560UxujKIg0+dDQm2/AQjXul310u+rvJKfsRDMmpOo0uFZ
xRhVy4ib3Ex/VnpuNQjlNHfOrHwx4SXHJiI07TsJWXn+cvZDMocWHH/3V7sTsGNoSQm23mhdRD8m
iAv39Eaz0YBzrmkm4UICBlm85QiZUDoQbb/quEFDB3H6MqLctWDRSCI9cLq+XAex3q4EA9pq8T5B
IqfH+2YZ4xU33Rc5SM0p0cQJpaQuhUrd9F9W/WDRPl+NNgovdZqcdQQN2rpT/HRRf4pz0XY/jH5J
fz8C80i4cJOc44lqQRnNVDzDYIhBz5qr2YnmDA3IPgIugH00QwB41td6G/GM5+M7jgqzSa1Bskkn
/xJPp4dtDiwDsPrOvExMBxi3xzLuD9vgt9d6x99G7mcULSa3Vw6jXfsvbvF/GC76mmAo2y/+wNR+
jDdVe7iGk2LCAI0gTo0IdW/W0HAyos8KPAoQevHXYHnZrLxUxs/aZI99jmxDFINswAYfIw0Wm16H
w11Rmvhg4OP5HBCbUZ/9kWb/XTpHluAX1zAo+M7GSTHWDwIv4Mb0NgUjJfxCXK2MBa4e0ol216zQ
T7+aBQ0MU3gbdQKQFu3ysaIVm1Ue5Vh5YMKi9jQc2rEUMzLe5jbkNFeMDj9H7Pdms7EOxjdeVfdI
VwKc+qruIrTIGbp6xznB9RHrai2dnIKDAwNURwD87f3FVELPq3+gMkkC+mzIc1xyPiXY1pH/76fz
yuYoScMm9G+kku/T/SJokdxQ0BpvLz8buPAl6yHinHN++bK57dYI52Uk6/NHVk+wU52BcM2u7aDI
SZJAxVmJql2LoGmdC0vcBaPR2icbFVz03TLFNZ4CREsSj90XYzj8YR49t4SbTThiQAmObUU85l3u
hV/r/Kowy9EVXkjVuDnl0HUzZ5IFbf105kIQO3DTjXM245sBYWTNe2ZqZCeAJ9fVOT2JtBfZW6pY
69sYuniN9k9MVDppC19vvyUrbpR/KISk8WvObfERdRPLHgCKnPjNQUQLyIMhNoHAbJP0YVokN6Qo
DTn+V7AXbRv7HfTcgPnXwmjE8+sa/fW7ASzsbICwKOcZviPdlcyFhuX4vBJ7ZUkQwvESCc8tQTcj
BMZT9kKudC1kqNK9HwbPYtgJWLOSjXX1hvhOby/mhfy4iyL9VpZCIFYkdlG3ocjSZqncukRu653w
9HHKI+xvJAhgdl/1A3bqQL16BNImbZq1B/IAlc4SaT+1CPjG7hNsQkzTBKAhYJmtmx4rHfpyiZ80
KVgYkwYCLoY330xL05GA32wYqvPdaE33wMrGGls8mzMCPn/R0PCgW1+U0d5BHlYIcViotNxOup/s
/bIca7tLNCqCC6GWVaAku2n3msRxJ7+6HfmXIU8YWIKsGlBrGbsQodQwxP675Addt1SxzQqvcE23
BMOF+H0xwa5dlNz4+RwAwSi+xi3jL65Pg8YlV8vDbW1KgPy7yD04DaFQTa40D/cjxbOE4sPaVest
p3ggsN3acyPBdGoPBum5ldToWBiTKCl0sz4PnGOXOtFtbjlqH4Eksemb6D/UBoZc03I9yP6jZyoi
B/MI47MjcoTJtV6Q4OGyLjAefGfuPXw8B7rIHVXVsde7rRGonvQsyWnK7+OvIOtQhW2PHuB3o6ct
ZB0ahE7419vbWiDnW4LmIo03AI7lLmIPfpmE9LiYEnaxKJ26bfo02l0wOyigUyo34Qx2IhkDSYRE
6hGI9RzxgkSS3Ey305U3id7uOiLk852YV+P5yFg3x/ZQzizXFyS++5CUABeUosb3hzPTzvgxdJ0c
LK8lQbmCfsXV8gL1RFbfMNiYjA5giJZfD4uCI+xKt8YiFc0AYPB6gmvgdjuKF61jalMn+yfeTo7A
xONholEKFPYhWCSjgzt5AdhQOc0Y7ba+2qN3kYAGcmv9sJV3WHBNZckcRgleMHavHPF5aOWQNFAB
bBkNz3KKV8OBNIR/sjsxoga0o3arrL4n1OouKthJ52O6IWyd2kxTFbDI3o2SjpkSNjR0p8ydQEMn
RTcK62VLizvLjEOmbOT8MG5RVIQReOpfYqHy1cWksIYicA45jGWvJUOxsHWtUMtoqOaiAUzhTuJb
4zTPillrFSQELUikRNVIbagy8qTRmGM6DUHrte4cyNV9ABKD9COf/fvRr1a6MKAcGOvIulGA90fS
fdZMTw+kKVdBtZInfigHgNLRpalzGs74k5b5HXJjJbWzXbYOfJXa1QbOoKTa+Bi9/Qd1Ij3tEtuF
OHyu582XIOq/U6Vn79365lkY2I83N6uLe3xyL9YEfoQJabPQ+qX/OvA03jiABcqsQYMQFBq0vvwf
FMC0GmTiHPzhAgSSEQ2H+epslLQtVcprOkikhLd3gfZY5lo9OcjyRG0NI2L6qqVMSmeT5iM8BlXh
bFIDvZJH8wbUverB6SiLcg76/h1ZCINZRD9lNFhDvtShjygfGVYZ5KFnQiN0TJBYrF9M+Bk6REQh
N/tIkmD4tFNkUBfaeMh5qtLo4yVOOqp5A0gQu6jI+rw9y0fmz/w5DuQPTwORK8GSbfxPpyom+gZ8
VgUcQ2F2GajY2cBDTAsINkyyzu6wQ7BZRXg25ftvSh2w9fS+JIaqzU+jz4JdfQBcuBBpA0UG9jSg
AapJhH6PxzvEpEZeg1uwtBz3o4mUQMeLI1jRvHV5k/g79k4VDvoUbEe/Nv3764V1nji28iKALBLQ
56gYNpy1qnBpVkv/FlpfdSHvfNKJBYEySiBNecrwXzttnq66ApIdOWmDFTxvDJULjDBrLdueaV8D
DlymqnYez9smW7/p7NECBsQUXvKQluVGQxHeNy8oHQ3mNHTG77wzo/iBSbGkEfvmYfihw4vTGUs1
oEwqY8Mf0sqT4DBeyCuwydINiuT7ofsZqESsMFB8b0apn4m0s2HxEZwhxPfGRKka8qxixAksagfW
Yh04m7LML50RD7ww/SCn+3MPnv4HVfUT1MFVYh8iWw6Dwd0tH+SLFxyw8wf9HxA3V2NBrVO5mobj
iCaMgzQ0W3RJlXPE3ANFGKlun/s2Zu3Vcb/guTj8yKAaB8zQLwkmdiniyq4nSxU9npsaq25euzlf
Z9m/20x4IM8wzzfwb2YOO7QSC8lZeyDRrrPEdvMYvg/FyUdOie8DxwUzQhKcf1xUO5330DIPq9Gq
TfOyItmXDnKS6onSpi8xh/CNmEMpjesM6nZD5PMmxB8h6tYewDUcn/DPg4lUEsUNDDHXODDHu/X4
8lvlt0rJ3Bk0Ho1RPz+5vV7QENzQeqe1LMpNtHkNr2erwKtjSDTiIAgNU2CkoF6/mpyMa3fXwxrb
x/nJYPqZLDtOwvDCXT7vU6EbdlYOV5b9YeB2ZjszCeXb7NNf8THc6KC4QF6CUAhMetESwvSHGjRx
6eJ9ZZNypXjYphIH/4ttZKSuvDIxqvAoD15MtgyqVcBIEnk121po/mGLu8Qc2hoPOA5bbXQhPBoA
EeN8yvQyVn7QTG1RS8wSqTb/x76nGvj6VwXNPFx9MximON9MLonZBQAyHSalmi+37SWJR5tT6RMf
tTZhLqFEhRle8iSOYMDRK6MzpJUfIHqv0m6C4LjLfmGzinyZ8CD7i7CLPuEG2yNgIFMynLSh/zzr
B9p33HUxYAHoQq869neBkyQaK+wJAuNd1JgH6ebNaHbe5wSBMpUtB6xlbI5mVTgVDm5s/wGIJrWZ
c7lKg6rU/5oOVeYvsQFvJVqAzJ7eDewIqa9rq6cndHT5/u74Mp8bdvrInppH5TY76nKQKQYlAQEg
8lB4PhbHNOPD/dJNd2QUlCUI6trEYmEL6AYkB8A2MydwTGq7PGMgAykNX0kHtm8clkzbybtW2EWP
xLgbrqm/tGy7x2Xd6o3j2WTp/rTH+wnXFSJRXG+hS8PIcGGqAppMESTbaOi/gvwJUXJ+hHTEHEpt
HjO3bReou18NwS7hUIrE7cJBiKY7EBFHdYioLmMcCHi/N0vwmSSvBzwpDcmC7JMAwuXYdtewocbr
wQ9LfJ9lPbMCABnLZ+i+b2Ulap9ARSU3msR3wBL5+Z7QnSOPUIHDtTa7vl3HoNeU68htPumfhR3m
Ak22imR7uUei8bs45LbM0KsxtnF0+0WcJpRoij+hmELKB0fcGpo6lLEHQuQeflwms669Au5xo+7V
Fqd9QYAShAyGD3VqgPcrqpGQ3BEkqGNJapCahlBO2LEdXJ/NgRXzgjfvjRQY6x26b13wixWthBTj
X3PI32rhLAzNyY8UNt0THxdikg8hAMzQSvrS0tlehSHnPXZnDB2ktg6Ii2GNuQHUWJ0ZsODis3Il
WcgiHWKkuVQ0Ja2RzraOT7EYn9EN8MXN1yXj/O/Yts2P/LBUMsNimUaYFoilukEi4Gpimmk8pRpu
g5iEEuO6zLvq7u5qcT+Riwu2TB2Qcu4C3MZJUQA6ewgWjGdlVzlibypS+g6ezeReS//X6XyjVzLZ
5Tu8xAl+o4gusktbVZULgp/dOnhzJZ31NWb6c30LjFqWrIA337mBRMWQg9bmvdJuecPqgiv4KSM5
g/rsvzretn9Il+vhbeYlG+LA/pzpdkj5YDX2RKob940bapRi+mmsTMKv60wHef/K8fo8gbGhEkRH
SuduPQaDxMRp5/rLn9+fKF4tvzrqmBqNz8xlf7E0xIlRcKGiev7SLPhomgDDwKJJARx/TYnbQAHs
IAm7c1wsMuIz5I0AsOj7Qi8Ry88DJdmty9BL49QqQYa3DkQZsnuUA2V5Xweghu52VHRmWs9smOpv
fm6T4zD6Qkje7bdcCbe47hx4SuVd/fRZETcAMPQM/48E5PVZ3j0JnVcyurV0PdBQVQwKY4o7855u
4TsMOuRHwRdbCtPnDeDw26ZI1e+4heA78TtfwIcmx5qH2lxCfiM4jIc+Y5i2zmnf69G6oyZlTSwS
8pPCBHljVxLYFG2TKUihIEtFEG5BCdTCC8PQxRPyPVIpBwnXizRGP/meGz0jEB5LuHfeG2FI/Orx
w2tZXUYJDW/hdGhovSSjar+uD+ZfJLJ48cmgdAbUCoA/oY7l07DNI8CxfSwZ2nQGochPf/nZRHqj
dhriEZBTZyzZxyNwBHZhFkZZnmPgw6lhQJyEDtSYncTsGONsQg5PtvWxvLrZTAHhJ9RE29sZVmK2
vTOkYRMU/VJMBVFjHjtMJOoPCN6HvogolpHszxieWOTFmATpm0U+DRynkzTTuthbOVlFC2IaVKt6
UYVgB5l/GCO0YDLKprd+tEwQqTNEcqdgs29TkTNwCZB1vUH2DpOW56LsUcWdnL+ibNKPTEiXvLDM
SZ8NCZo0n8MxKmgzv9qTt6pqonD4aMW7r1zVjYZ9fuC6acoux/GNlpSMHONmf+EN+fr+ex75LVTn
yx4d4qQMXycUHpJWFEyp1NweQufARHkHeKl1D1CTrjL4g9x20TUlnQokVy85TLaPgm5vAaEldMOi
IentwreTJ9P768wLRJD+yw2R99KI7Dfi/3ibmcGgpFmLqtVBpKnNkK8rgvsb1KAmgO9ZVxDF8IV4
q+mlW0xlb48doSQ1HtzND/MSxQuQGSd29ja14+C3R9hN7F9s3h4m4uMX88VK+nWKlSVdFDdvqTjP
O/EtVXlARcBcD5ndLapcVGtpZ49c4C9dV3qn8QDR+bPHVPUeBxxtH6HUKtUz8hb4RColqnWwHF9d
hPdLVGOE791cBaN5We/bX46T80HwQ99CPdQCcR720xcekdWiFNSlwVk83UWAGeXwlNndDBYWYSBm
cXsbqUYJk5TWw+WmlcGSTWsJtUpeqGWfNcGIz0wjuygl9q8iPYo+UItTqiyhebaGThF2iEQ/mxe0
T536DPjAceMP1q8P19I/m0nZSkGhvvvNRwhCeplmsQ0bTxm3L/6leZ24fIFNicGqxI8/f9b4DUY8
fqXVqE75umTJMNaxi9SyYBQgYWRs0mIwBRcZG45nrWJzD740MYgOjugLowLrXcZFB+jFyVu1yvc/
bEa0VqaEt46gMmoAfm8PnZkq6CRORrmip+GqV+7ot4IXTPMc0s0O5fYuiI4CfEcZKgjakKdK9AlY
ICfcTOgbe4XuQ0uojVU4BBWlIXToa/d0MDwIS4AcV/PVK3M/3EHh1bNp/MwglOonSLPNiZRTZv8E
PfU+GklMYd9NBygV6z4fcQTxg2XTrMomhiJ1ZABQHiF/3oZBsBbxwx7nh2aanMU5knRQmD6lCour
s6wOUJ9Rug49e+Vup4E5z2WzoB4wS61x4YVK9SRleuRhQ662xIO7E09a1kOcFzPHUByPNJt1n5+x
zisdWaiaqAdjQv4L9Vr84/xkjv3nvQKxWh6CdgimAHrYjnEMtk9AWClEfJxjLKMWIG+2+DR1QgAg
+TIMlQemXSYgBNVeaaD46k/5Ds9xRiATxSy33OZdEEB7HhKudW2C0usqJVT1bAaTSlZ+RyHRGJpY
2BtDhMKuD8zrPvc/vtzMd9sWJSDcZ8f1yLr+k4+UVz/Ep3H7UEpaTzcFjc4dU+vlzBbQ2Al4ISBy
u17XtxD7peZv6kNZ3/MHumrSLujaEWOUy1lrchd3VkaK9AyTFUeyjeidPaY16XG9Nu9V+bRLaHow
ZmdA5ZL38QXTbudz+EDtn6bXhnuIpdNPfudaY1a1AD8DJ3ZxpWodZ+HQgEpQcVQ/xO9X2YnRkR1K
eL6SlvqEMVEtmBQLx4ELxVlPOAseiAI6P+26xL9kW4yK2weqlXIpcpQnK2UG8s0F0Vqw3Bh5Rv9b
HmAevj3ex/G6aS0rT/BDtu553XEbV2OcI1rhFgNclSG3EvwqdIiHv0quYyWUMu8HLzFy0EgKILGB
18VlIniwc5I16aB4QmhP3sgctKuDQZCsusSP1amDWL5gLCRKXabT1c/7izHTnioxKOcHV24Fpn7n
wE9Z5C28H4MZg3jQq9y3qzzmk+jw5f/IM2QF5lkkwfDld2/+HSvxaT0D6iBeu04i7EiqIl3mMK96
LtMDWgIE1IpNet6WctNnHyk5X5SOdsdKK3bwYiqtqJ+Lo2hH5kJpNkPuweJEKellMDfBgDYfGGZy
6wyVU13MRKb2hEGLkBVTm1fzfGczAxhwtMwyT+vfr1h2ez6PIET1wujdAoWerDCeKRchN//d/M5a
PYTl7K9+zBCnqXfnRT5Voau9SOEGKkJck/pWwFwwRrWBIbGPEUFOMWvrFb1tYIE+QfYtqpg4KGZa
pR4vSUiKak8ixh9A2PTK3kUD3CTIuUWd88jEpfKkRamc7drSJiIGEEDULdQo9Z5wXDh/Jkg7DgDt
h2icTH9K/dIPOsnq9uurl1gpwSyBb0nCkuOjGtkuyPOUYQ07k5xQTHgcPoIbajXKZ5btum30fsSO
NFzLGGwcjUKeDmgG4UfA99KIRqvfS371e3x/daPutsYSgG5n3ZjT2HRFiSWHKWxAmXp3+4K3M5RE
8mM2uLpLGjnN3o3JYyy8UA3AD6H2QlC8t/Pl2k8iuhP34m2Zf0sH3s7WmUb7AYVdGAvO93QKCBEX
frF4fG77i4KtIcy953pCc1sastV3vz/J1107g9otBOo+so0MwApOAwOUMWRn3eGy6PK2BSl8DHNV
WaCHWz6K9uLjT7bvIBbUl5T03RfyibldiW3FDlmRTIr1Qv5QnzVMOagelm04wAZEvuq04mBL1Tdb
W9VDZFMt5kFUnXNBkAmrdWEXPfg1lSdQ5It5O1XkcQgiTzbD2CZrbWXDqdcVS413VSDMJaYXV2sV
EE/pFAAaFq15s+pzUpgj7ytmB3ImXIpg5XR+akZ8f+EyQx+QwLQnr2LWyxcUCrCCsp/E/Ll/OTL8
eZw2UxuvmYVFhFN5aUIY0+l2dzegHrcBRIW/RMyxu6NlixpNerzvTnrO3t0DdpmHZPCxHpCaufVq
ECEAeovLRJt285R/soDu5c/6MG2cRc1zmG1ZQs6GRAdeoiGH7fywDN4YilL/Ur6cpNXbjaBoo6dy
muoek7byPnxqE8HafOxx+ljBba0OQae4friySfXseL9yHsXQmBFywP0JUecOKn4vKMA20Oz+eSdA
+MNm70f85uadnhN/ynjz0m0JpwBl3TcJvHLuAWXYj9oWhbkxthkiccGln6FVJO3hoHhWcgTyEvhx
REmIjlwBYfVqH5XBK+TgFVHo6fRom5ckgxLzT31jqM4003Lgk8qo9IsYPsXq7gA5ZnkfthUFO91J
pEYh5KRg2LvMgKuu7hG+EvmQEt7hU0+oy50z/V2jrCDMSXpKYx7kD8MnFR2376DjwnuaBn4MMToD
Tg5ZUi3KOrySDxJxmQRTtNd3JefcYB/pvEx6VhXdMOE0uXOAoOLhYvzrDWj67y+4WXB5JWdmKF56
p4uwqOXHt/5ZUCKX+3+8FPsKZ78HcDzLke7oOhYxJFrGaeUmwPxurjAAVKKdafM5r0jI63sRaLMn
Tf6rXX0d0KVOKNHsrBosaxNznHJZKDVXRtFIOKaxJc0JRuaWi6xUFDCJb3uMFCSMk59HVaiW3vKf
A5lwke33WmKLF3iv3rRrmcj4a8HnpSaHLWkF+Bty+vzVqlfLURjGb7ze19UACUqJJSreLZ2itiBV
KzaFuCZVfmwjSHx5rwqRbTHwjRnF6tBR14kwfNlptCoYjr/zd9qd1k9pcFTTjzzXf9RRdolquzYB
xFXI3idD+cPMLPZ7LYsMneQMbsp8TO8LRkXrYviOoe9V/D3MjU7nrmOYKBPAMTj6l3wxsJbuf1V4
cQtF8GxnhMLqrkg5y4AzaBlIlyGj9TRGGxUw5npSkz9EGLRlJBgRsK0gLyG3XY9TpUD4z66L/x3d
or1yaFqSHFcMzPsXChq5aMwekgGC7RsXQ1OXv32PC/9EHXYEk0ODZODy2lvygHguS74GU6zjcmwi
lAPNFT5IIoYxRJqVuPWmntgkyj/TxRSzqCYn6EGs6Q6crGXsAJfD8JFatqqDN8yQ0YByObyJ6aKj
GqBuwDgoinko0QUTc2+hRlNvGrWzZ38VqLx7OVU8zzco4sa5MyBCRzSwkjtAUXYPOL8Al3cwDMIc
q2GHRlyaGDEQwMqCHm00VsX9WhREFdYVOx4Fub1cpHDoe23ckfGuJ/zb4B4picaxOEmwS5pmJn/r
qANEP3JAdY+mbsX/DVv3Y/8Gz46uNSvFGY3oN7f17i/3uuyJb6V6aRjGT9ZUBxPQAHEQ01FcEmme
OY4+dz7iO20O0xnY3WIja+cAlpqo7sUTxY+/TqF+TApPLx7aaAvRx5iBg9IuoL4zAoewrpHkcBqC
27q6wbyowERrPhCu1t2W3oy7nZS7EJpbXcUUHvZRPelbe43UA8yF7JpaFQDkMFIt2OSlsnMKziFl
x49RXakx2xYSWHuRPCN9esukfnv1f8C/eg3JJ3TR93qYKoxLi+d1JD5pGwD/tHvsJd8SNxliU9Tt
n+vUW5N9JiSlb1XEP4d5gzIiHCvLN4151/jVKP9W/fPjZBCQYdeZ+JfeXMukKb9pieWwk3Maoi9T
gaqwGJg/OxI5/RoIS4y+Glezw+MfZ4MPsdgVAoqc5OeU7qRMVGDTcV7dnyrvksyftJrkRdRw+iTZ
Sj8zyqJDTESXgSwDTKMMjjRDH+chT/7VKKXkB+vRTV6ZJgL5Y1zjiF+Q/Fy0oEbpkrKHKBZ+iyc4
9h7wDW9jPzoy4ZKi7mFPe0/7+jvm7/KdQEfFTgEiYT6K3GKdcp+luEsljtERsqjh5lZpFvra4QZi
8pWx4NGlCGNIIP1rkiZDwxMaof4RSZM6YiQDEWVXqFmW5v115Q9y8DtMdXnq7gDWYfjx65L+yo18
Uu29sByaIGc5C2KP4+UtXPKjAyLufGxyth3SNk2lHPNAI/mA1YFRXW4ro3T8vol9g9ob/Dq5KfIY
vQZBlX6QXVpfOxrK/miHN13wx7wvX2P8Q8+ENby9h4U0ErpgEVJvSH/q12lQDiE0m35+AoIQrZYb
zBx/qU22fff3v8xP5JsDpoNir+5R2njowpVvFJsm9q/tV1Tbn+5sRGV4x4xDlfDx7NJWCxSw94qD
SzaDOUAKzXyHyvlYvoAO8ENTgIMkobYfIdbphP9hmD8zNY+HUgKIqcfQVEu02rGnkXNz2cg/qrgn
FprVlw9+MT586unsb8sQyMHfKRynNWaByBqdWNhra9vboEl49Bn+2+99B6tmPVVrRlym5+qbwE0T
TyIQHHwjWzjwt67tO3HTZ7VxCQEYz4y4wrUzzdUrR0w+nbIz0w93Ii9qxcO9UqCLYlYPJU9qV2fN
SASOlu4cP5bZAFcYvjht8DAEw+UcdsuH5mL4GUY6X9kh5nvFruksITaWDy2XAipDjgRqCpDkTmYW
BROe2ecWv+fJflDwka9rFHFDn8leeNYPKqtsVfDaAp0Qs1/3dS0y4FVYHM5tWWiyCeNbyhaM4M2c
b6Jl03XPI5gf3MArjYy441z1CnP0fgPDlgeMQC3jaelHCzt2KGknHt6UvptuBM0mnwnh8Dr/wLjB
zX8MIx5ujfhfUwDdsuaDTSaVzpzpmlCjrgSz9X2iBUotsj+HnkrEIDU5FjgF5wIr6yM8zcfXbKcr
9R07b40aiAAWR/kHRmqbtGgFHQsa2b9pb+J5zDdk+mraEr/R+ARHe6H39uqUs38s8kT1+5nKeBAf
EnoMvlB8/iTeF5IPEoE1tiPNJ8Mg3wGjA4TuttP9rb2AbRGaXLM5i9bXB95nuXQNiGZ/6giJO4Eh
3/aRq02cREIoQs+OdMuzQFOvFkKb2R82g7+qs56YX9JGzGhFooZXx42PBUFbVhQ/TPUKw28TFiP/
2Bw28x2HY4KsHkeVKx7rHYxBCNnOK6NeNqFEJJsGejYS5XciRxevqs6yOLBB+3SKd2lZQb50HzMj
xSHlO93O5TVRcI8GcEapMpu3fBbN2EkxZrB6SN/MuHiBsFV7zgO4iEsVRJGEluxTM3E9GOYBc47t
uHIKKEQ54tDt7INPnWvovnEi7z5hYcbSQ6GK9uc0LxP6amLmPcc9NMXm9IMCKt2U5m8B8rz41KmM
NCZg0tEdj6y+iH9imqTvADsHiaHx4lBHShdanHTtANgyaCoktOHNBPJfVVqbNK36Xo2zmFWDY7Wh
p0xxt9xlgLG1rYqRaq0gdmtaor61iARwhJ5BKFPgZTWg0c2lB6Xo8FFHaiuAdVdubFzTmLSMawHl
Wrnu53/HgDiyxSjpj1/D7w2oQ2a2RRlXmihfQuLYE9K7s32pp3KtN1nCDJSrXV9dtTNa0088no8P
L8OM3000yaJP4LA5/XR8ApxUl+0+81xJjHZcP6hjU1ofoZIcfG33B4quzeUyl9IUwD10+o9kbRkJ
wvlAkAjUFCX1v7Ymg4ktmgforxlKnYfs7mvqJZFRhRMHEySMCzFO9xEWKhRS+crQVLsesC5uGfV7
VoQkM7JDVlbQ+R6iQtyoG5QZw7wYzXG2urygeJTSePYfh9O8cVAk/ZbWzsTLYkKGxM2z8X6gJ9AE
864yK4S4lRdzhdETMUIoI2O1kGF39eNDNqR0FxVWHYtMpFrO7L+gRRM+PrznnqECQLvYbCc+qCH5
XeUsIB+X3QB9EdNDORE/GYbDFxpObwU+LAcDuZfYMqEDtx7jcah+OEgjClTNokRQ7wiswzsUcmEg
73aYbWUzH95DcqCbYgX1OM4YOZQnE0henyL/0K2D6BqP3+/E5LU3kIXb9E0xp076o5ggpEKJPmS5
OYeEV5bX4Pvw1g4UJ4dyipoEWiRHAlJLZB7MeCuNEb+llAu2ttN6sHvXbX6aVm/1bzb//s+rNPo8
Skvly33152JSKxUtxoYg1vuggbhqliDwxGXyR9GVyK5xIur00i2vm13Lkb0RAwCMrsYT0a+paTvk
t/t6Kj+c6N5mmmXwjaA/M5NPuqTOzayTTezzftpFOizqbzatLu7hPhtoc736MjYfv8pn3TdTynI7
y5RERo7HGttPwVxf3XPXySypRN+tmtUr8+a1SEEj2tUuLYgc8T+0HEZNpWl7tmKwMlwIl2GIK2vw
NApsXNVTfsR8gJ2Rj5PlcBst3TWJLZCRjIS9uvR523w8EhnJwfVwYIsBJYpQlnKEj5CvBB18bpfD
BfIEzvEArRuGnbRbewVUyaGmCmPNd5DeHIRRBK7aIwQcgSCo1vXamTa3czCYfWdu7fsNs0UgsI5W
OoOrW/0isJWGS7CSbs8BJ72GQ3Xh1yZEUyfzj1WnQzcWzMMWDMTMXZsO/FtnAOJZlILFQMbzL/XU
963gYw/KM70y1JICDuBwdJb1/xMSG8lrJVx55Nz7j68NmMexe6ba1NpOI7D0JKT4Zejf+pGMZOml
G5gRE0jCxkUL8X/2vw2MqDgD5zQqN5MQVsVbWgWdk9s6Sff/DRv7/HJQ0ZfaD/Gfd0fV7yR+cW2W
dBBbdYFbNyLVuaD72UCjQGseWyncAryHjtdoQMpdswKLidkttBeqLLW2xhy97H1gSB32uC8sr/+F
txXBwqivukdmPeoXmvrBlr+J+nw/n6EKYjmDXfJApbzIkdbZcHyn4MM2IjL877K3n6gHMIrLa9s/
68F7pd5zW1mIVLMz4BseqV6kDATQ1W2aIEk1RhgZWvvVSxAmI60XS9sso7H8r1sz1LuVKyNais86
XRcWqjez4lBBBEJ75ARNX/wm4ZgFT02SmHdl2hNbhlRDsnQ4LiO1f/hY0A5BbIVRu6hWxv30M8iT
DmW7GrQ1MkV27Dkfon41U9cENO67nvY3X8wRa7CzkAku16oir+emosUanNJMHEQUD0tz1/4wooMR
O0y8qclj3nyW30RQrP/qYYlfv4FO527aW7txzuqq3ySPAg5Vi25VyXfEM6uc3eaJxGUyKmetV3u9
ylby3Bn99hOOjavw+X1sFmp/OvMyQrIBhhHhkhht1UOynrzONKuC9xwf35fH7Vlb9SPXvAOeYqUh
wf9tf0XBrTUpVDgu2idHe3wLOc9QBrJ2f2tOyWhTntbH3Tsd8Py8+j6i97HS5c01oHMw2Hssn2TQ
yOHKCtrRCknp53JZQ7jIlFmhS4rK7JiqDb66tHQQLOMrDUiGMkHeTum3PjhOpuWDT1oO/+VU/hZG
NrMslN+ali5+b8rYD9B//dXUp+ewQ+NX2oxljWvoUZ339/otD31tjLuKXme+zJmyjb1Y+teguvnK
Gg40s8ru5GejW84+wUbCSbiG4aOH9FfpyZRS5BaZl++eGf+aNObUvmrftoiXZXdtqriDm4qzs0k9
xI56BJlDWlYQ6DLdJgzAb27eg7mXgI+2os1yjrAEsDNE447/lHAjI5iJhX+oOSHMbbs7FTjtzDrL
ttNdoVBbhiv95Dmsof2gKaJgxBoMWJumqI6h0GCvn+Dlmt9muCAfGoakb6sUEToHELlylF0Vb2aD
dtq3IAHjNjVSWEhJlrjTIz5n8PniT+cLcucUkzZHzZiP6AFw8li4COecfRsuHcdt12SYrjkYS0ud
qToICGbU0s7uG+8tSz/ZQ3YUZ6fUueLvI6LTbmS9QLtZyq+LodZrl1CT3XXnfAURlGtSTrLT06hW
U6At8bPeYSJ8koC9/I8WKOm7VY81hLwfLIyfeWdcQSYpiHoT8sNAUUFXvGUXzd7uHbMMsuXoeASL
+IJ2uZGvOLk7nt0AqBIYXWxwUZludaUtS2TUyRUKd+Y93mFqc3vtusewguIzD9Q4xHRe864X3dx1
HTqmhZE2KCL0Uav/hVgIkaHtX1rLVYJudVxYkn7piZ+soqX9d+PEtvQUB/o+2AqAWCnfJZTGWIXV
MrxVVjvU9KlEKwRwAWEqzQNVXqBfla1OUFUvFKO9PpqXvzzoayVjLEDCFzfAlR1QKmwNkD3SXfg8
aQWx1N/CsAKbEt2YEUuUP6u+nlwl2+/ijFTT0wDI+Cu+Sh6OOmLphWnxTrE0MhdnzYglyd7lRRPT
KF2lJkOhM8efZWM0Qzz9QXyVxMP9UPcsZm+7V+WOkXQ9zy91DNrGmV/NgxEkzDSWzX44Za4/atDX
0uzSekq8vkEeYOTLXkbhri490bcpfAgOvH17gu/+AV1cvUThCnauPoreCwsAhvcfbwm1Dt9zrWBZ
/7PhVGCMJyT+pxxcioN6Ws7HPwC8adkrGgpFhhbMfuNueEgekT+0nnqva5IObmvcT0yEoqFG6jYV
pR9uKHUMQeWZKIWDugKbQ08JhywMzJv49jrDydB0UiMqYpLY3xN48/2zTA+ikiAMlLBYWkt2r4mH
UYA6wI4j375ba73EXQGN+mcyiuhvbDjuAvAG8KL0HBPpW07xfeCu1bc3YYucGbXOlyJSFSF1dqnz
xwASe2zxQXJkMbxUyp6wYNXlo8mI3Y+dNHCMemBxq099rDPfrEFXJ7VxCStnHCK198oN4IZW32O/
wcJaHJ2EwY0S3VcB0a9GIjhztR3HSkgxoqLCT7tBgMwxkNeC5JlYYENqZZtwYaTnafxVa2k0zFGH
J6I8/Q1EdD6mUCPzzL2Ly7eQY0oyXiaapmee1EdIGLAKAxEwUJUEudsdfJAQKyCT7HqAKleGOK6U
9EAEl+gYtvevZGKa1Ee9HwaXZvaZDXo6VT9z1Kw81jv62ePkYHJX+kEULmjA0fLwmATY2q70S034
nmDZDF1N9jAP1AZyLAO7jqkliFMupr8k8ByXa5AbWn9rkkZaQ9578Mefu1n+q74a7J/9HamuiyXw
/10h00rzfW6a8ngxSTD66HbX12eEye06w6lgBVEBHEuZtDMj1ZEkzUmKWuEoVSYSNmeLw70Yadzq
F0/rzrHtXv5F/x/SJjKXN++nurLEd/qYyWLLa+uo4xUL/sxj/uvHLMp0PsMxveXz9HiTDxe1Pq52
RoDTC+eMn5bsC+CUHImwF2AQgro+qxfc+CXQcbOrm/M4cCL40yh8WH+8ImYJvGNHwAWus3JuYbXY
H6nzdcNUG9xOHn6XuzDZC/SFwBmUnhJq7KrzlTSLf5VSXF+6NnTCVqSrXqLCDv1svYq5azY1PLir
KbRYsJDrelIA2JLwHQuigUjNHZCPeTcVHWntZAYu6bTjBqqY43imgWhqaO5lm2l++1tozKkKtg60
7x/O+jE/aYvNyU8UkeMOmMrLN+doeWehm6kxJhy/Q3Lz2I/8tA7zO065r1c77GdL1kIgy7r4jeZS
Umm1Ae7nm5IvR/wB4FV/X1tXJjV4tIcz3D2q9sKgcn9o2TnoXBjeB89vpiti/NqqH19V6phIP5o3
qYnp7MUbIjIruM4nNC+9UyfNbDIgJt23+RWKTmH/p4ZS5WJjTQW6Zmr+bwlVBokwCpy7WdYSCBXL
SMcHyAXYZ1mFrO8NGSl3O776Oxuy4ivfiwI9hROB9TtWuJapIi5+gpydM9SEIfLncW6oiwMcoqar
OiOHkjLzOfUYyR0k3/RrBmu+70rafrJ3EbMzoiEDPemdheN2W3xK387/QSgNvxnmerdhTap/qL5X
sEXCHjN/eOgcUC7ojTuNvDGQauxTpVE4anUoNf2hntKmAqhoRFDSFDv1ylaxSZNwzHO6hdrHktNX
m3P4eMIsHtzmbZiHFSlZIB+yrwJsx/t2eS3m8d9LKoh7nprOji/Zb5sjr+cLMJYfT4DvUJ9oHXyd
K0Nkgm2gCVlJpDbKPm4D69kVXXQFKLNKmTRN6RCiG1Ecy7/G0gxpWDgU6BWc3JPpiebm0iHi9zdD
+NSZNlUZD3QiPfcN255HKCjM2CD9jmQvlFX5onuksEMnq0rnAfhLygMe5WzFLZuC5z+/jlBZFtsw
R6JgJmubaEiSxHnKpsjZutwnpuMQx4ct+go2kvCDLEGS/aOFzAUkgqweTazy8/UyF1Bx+BKASvfH
WIAwPx1SNhsIxjzOjgh/lvZ+zjEQCVG5ksEFOYPFr6fKh1JGRnMdfPG64HwhjrAI/w4RInEgBT/M
jZrej5vcPS8c75H/3l7+cRAR+vsCK17w8NS8TSK4p1r6Orw8PRaA/BCU6DS5nIfN6GWwJWeendNs
ZdqddXRPzysOj3XjV+bJrL+PkwvySxauInXk0FL12IiTzGf/PxCGGT3TcGGKG5LMj76cwKdQPDcf
1VSqRnh+CUnsfVrmjGz1sp/Huw9+xuwlvUbxT2q5DJL6rzK92gSAdtwXbhaemiqM6ZmmuNSb5Lut
iHdQISqB2f6krdsDr1NITd2W1Zi+xIEEN8Ph7zrPxaFInwsG5RXxChQ+vLKBylS4tiy66SIJ0jDP
cLsA1I6b0Bg4KdmHP6oOwGBmJO2rI0GYpcxnSKvEuEedkCbfLpkURypbx7rpn6HTOdE6fEHgVw2J
2uIoWiqEWhpbvSjHdEmGovT9xRZ3vKUMGgoTkDkJ/AIr78gpUNPOR4868MPg6XOe37qIGnvlz1zO
4563gp54qJC/otfE/JGavGWpx6HqpKGQ0I+WXpkkYkxGJfrC0X57gL++agaOVGwSuKt+ui74eGe5
XkCZsgxBRS63zOzQx9hC5UcqSboXEfsu19p3cf/0RNuPYHQXN07sCVk7HNXsgVskGBX3PD8Bc88S
mxRhoZzsIsOZs89Do+4bdUbJ37zVSCGik9MGHD0VEWPSDQePtP8+Ly/Keeljq1nNXJNz326ysb/b
Xv5ZQbJuOltqCEXrxRV6hkytaEx2sxlQ+Yq55ULm5thWjzz4ytLgUgY19zQkShtSQu/VGhWhjg7f
TbhKcYXMCh1oWiZ/tOXTrUk2lVRTnFuGSfDa13dhFqIUIHdI2JGAQSBhsWHfRFIapOVx0Ah6G4Vu
1Ny7EvAoDqg0VrGNpif1P1G2T1QOyGzIWW9JkwuDvEJug4d3YiqSg5yEqw//LG/KMMDFZ/xHt9Yf
EFelKtOZKGHsexyud9LRJLGvvjJS69qoIrYRh7qJ+uNiBReBIzAk9myMQMpCtMZ+kKP+gOmPoVYj
8GD0+ld5WuYpobroMyjop/XjtgvgL0eTlkQEFH5DHoI9ma4dwnxvTjzqXfRnJLgceI6oFMuoach7
gsVO8+ZZm+uYn+LeJHSUx1d6kr88YIe0y0Ja69kE5jn0rJ5/6Pbpp5xAStAr3ueUnO5h7xsKDMh/
6kpzL4h2nhPc6sI2e0AZSboaG/EacS9jdlUq+Zowk8FEbyz4dfq8MMidGddiZiThmhFvdXrfeMA9
MR+krEcyT2WLT0HqJ65kVnn5NimMdeGG9lE1QmOcaLEUDBhXslrzobKE5GPgZTCr+x4mI5aqdT8x
PP7Ohe/eZ04iKNQXSK6FBPgh4knAucYVTK+P/bGsRk/blWfDK2rfD1YjHn7idkL0qADbmwhUXl+v
H7BQ4dNKHitqvRob4Qo2ZhcUp1BLQjMF7f3k8zBEGiKzgCXoAnpRnvPgoBxKZyJ9/0aauvVyWBsa
5UPuBYofrPX9+UnYoa8+Oc1L6c3zmZn/y1hiv+KOTED73s05NStMfbrbXiYJdduoLPS2K3RoZF45
NW9DyPlj5nRPrniKeo/sY5FDE3LZTkB/IQYQKTbSs++bS6jD2Dvlbted4mcCxJSRc5Pqj3+mO8/p
AZ4z1Ib+wfHxRrYSwjOXTLfSuTkTBxoa2SCfmUlFWm+Vftz80/75hlGIjr+sNq44Qe3lXRgj3dsC
nN+S90w6Wk/Yj2Xahv/rVP/9X/K5OHvC8/8wvRLBMStFKuN9J8S8cbDhcvnPXbxdwx/AXsZ8jAqS
5qtODeIZQ4wiie7EBeP+c6SuvEsbhT3dRefEC8trFPC+qwTAvq6qAPjgzK5bcy+7SxblzkUm9pP/
RGLjA2mw1Xj2m0SpTQw01AtJuwtFMco2CVH7Zqf9v7+oJBCi5RlLWQsl8ZGiRG5xPCuX+0TIm4BT
8kCHlbZfReSClU+iGObQCwe2uhaIb1Ww3Dr6MMjMFsSeCj8DmhpDfbXcjthT/Lvx2oqaIZYnEADF
3Ozt4g2q7H0NAjlB6bvobPWq3QLF6H0KeoWvAJCQ1oxvQUf87IbyMaCigi4niayDApoHIq6D97Sa
KYkH3T2uFOpWZjU32q9vDPYp+BX6rhPc7kjXrXEqgaKm55ACYVP+PAzSaPccB9sjoi8hJo1TAra/
bgBmKxw0jgy5F3g5AQy+FsUyNIzK4afx/1yRGLiTVRzbgkGkOygLVGuK+ZZMjJFxETbnnj1+7ATA
F6Y9F/yIOJ3PGusst7pRndNEtzwXaBDO6NFtg+AKv+cJj5m+spkRTEQbdSvRfb7OXqrZtMFaIGEo
mS8OYCywihTpFe1BwCAT7RU20erfYrUlYYCmVYtyZLxArX8XvOEq7MWUZ3hPD3FXpJ+4D8o81jSr
D6U9Ukd/jhhJCJRy4dPYyXY1+8xg2JEo6Z9tECv64/dpi4ToUyP3D5ry5q60y2P/kDtPeQyGXDqR
zck2IDY9W4F2tl73bHfU3Ad9yXrYgrFUAfrKuIJXOPU9Ut7QRyWMePeSRAJUwCmeg/4uSjyMjBTO
tJpNKFy6s1iy0UdyuZS2/cstFCdV95mNOBu4QnPRFoOiyGll7Fx3cNvGXMYlTbZyN75C0aZW896I
B8MthNz3J9reVU1Xfhor9JWtYD9Fo0PCTKVvMUt2cUZTT1rkLcIZbTG0QNMB2ABb3MlQAwpken5i
VleEoRdelkSgP9fH/xs3C0huuEOEbHliOS0u7+MOQGEHMaVEtNDwG6aEl024Pewt2c3fDz/n6fzD
qwtWlplteY30E+YD1D8NEGNM3sh9y9tcmIIJ8v9ToEcjiuMeGsbGBzdi7pL51S0WVw6yw2iSimTE
EUj7sTVrDWGpmY0HoF5tNxzxGrLJ6/JdxvHFg5WivaYYmanPrViKuZjwT6MDjvPBMhYqPSzc283e
ABCyZ5E31J6aRSHZVqa3L3efVvHY5f9ug1oElzBpEMz+l80Rcr2/qGOIj+Ep93DrS0dwmGOzHsLw
qPDdeuIH4SpoqZdGh2o715X5vzjXHRjCsBH/FOcVAgw+WDisXrgu8DKeaaLZbz/MORMyqWq3Ovsp
dNnFgvLG+nq1pYyKIyOkZNTzyOYNJy0JfXUWh0TVnV8ql0Du/oDcvfDelCJ/jfQrLy9PWzUJqNkr
bheRZXJ9ReSUPPWpxNgWpxr6s8ukYy7wfll/8JIBRrbLTq1QyHaT98eI7LzxyGrv0Xse/IC3rhN+
bp+/XGnoj6yalLth3aaA7gmVMFUPxHh1kYmGQOBarZWHNDgKuqTJ4JACIRTBIeIdppK9QIt7MLVz
8gghp2XxuVshR1k6EXXWJl3Y/SMyP0/2NXmpoY2sUXlUo+5R7HucGwq3EHSVHEF08SUr7QFQVYHC
Th9PGjNJIlosbwlw3lswVE49yjehdKz3eUlYgCE1+zm+MORXw5DZkF9DAIOrYetoeNHnl9ynadGh
/s9fWMyAIr3zTFodBOYLexF1EzunW/BL8uOIXVPl9h//NpJKi6sT5HokfZOccyijP9DsiT2SaySp
hx6RL47pzsO8mkZoTzpYolDCXpjio4fg+SOpm96yLHN9u2OXIDVr3tL+Fq2RoqNrfdNSujN8PfZ/
jvVcAnJ6Hcby2z+GcKPa21Op2Gih2XNFJ7iTulMnrHabNjrMcXsS7FwtNy3a9z9jiQKsN7cPnqJA
sqQ8S+46v2kBZ84GyUvMP5ysfjQIPJEplFTqx5ofoNK5m3w1cqVy75f11QN4JpIFCe3LpGTRXNVI
2pzbNiyBNh25dO5ngGWfXsi0mkjlo+4N++51GaNNtKduvrR4WCl4yYO+kPc+ZDinWSehDveBjnKm
qzMp3NYUQk94u0+ChqPj8CWQoJWceuGtMWNY/rl1ojVywWb0w7jtQE9wj/lQjW4GW1twCpNxJrc4
ECvKtwyc8lNJdX+Hs0II2GtmIJJhkP5x5Y6Z1nnC9wpNJGQVuYggdCOSE0v4Og4lR5B3lFAWgIxl
8GqEI3DCdK/rL8V1g642FU9kX+CRT4IfY6Kf/mxx6ge7IvyFi4cM76H3AbEceWwWfSYJw2nFzkAD
G+B/0DnNRwMQMvy69rIVSumzPVgkJn9dgaGnBVsnt0xelanXR1DD0TWlHCy1hC5jLWEYRELhe1aZ
esL+1psTMooMZRHF7AGjC5yBIi5d/L5KRM9ECAxCAADP7NH4um2CLcQJ/O796JhPGgWrAdCGmcVH
JrvhaNTInxF5ccFH8DgdJXx3hzFKDbHEWAd9mxU8U+BU5O0KaAgC12nSWJeRZSzvRHbxgPxq5nRg
Xh5Pb4ZwWREN0tXzrIGrkF0o46rBcI3eSssfSLt2LXxTnuoeva0H+BLBDHu/bVdV4wGdV8hdWT7J
4PUfnsaOZXV36YFgY74Ta9ihrSPehsfX8Hwgt+Sc8lMJt/PCN9kz0y0Vf4rbO5RqTvsRnBObTIwR
RJt07vNNk0m74cvNIF2RvoUV5jkUKlUJd5LB8tbzh2ydB/4wyidknLk+rv0y/Sa6aXRRz7idL8k8
sYgS3JC28iksbpuMV+mkFxfFFLi+p8XeIMY6iSWAjFk/hkr+euPsBJA4rQenvZaagg9+mtDV7cJN
8StKPRQxXb6iZlQSpZBgRMWCpU2cvRgyI8thpW5xgRyfxGci9FXxLfaujl4YlfMViEtWi6hI02oD
ruqYBW59Bb4lmXoGuRkOmeIT4mon0+z2xRpcwtMSWM970XE3ra0zP+AfMyiRMUP+TsLJhgQ9pcrD
FJs/30xHNmgF9c76YQjKN2IM1WO8SMsxvP+ynavOuObVdT65Q3Iz/oB5/9wsOaLWwIP+4Cp7UAeR
5olFV/x6UeBxetWk81v+Vhn0Z+Hp0097aboW8ubQbeHqlXo9vVYIVzI+thg1kKQYuWc0J3pNX7Tb
e3ZR6B5faZO7spyWTBUE7Bg3gqtRVYzccYfi00113oPgQKWyzrytIIqWk9xmjjvGobNSX0i0ezh9
WtxjFEj6jiaJnqP49l+X4X1DzC8wCA1++AneZDJmlj0bLUCbbkdsFJtki0nnpPm06QrZj+YC43a1
jdgJBreX/OuqH8eU6CaXnJPVHGA1oshRluv0L5Kf2mVlxvQnYuvm9QfCpebU9aEYmFcIhUQBEMUk
HPvGSQUUsJjxSR6bMJXDqnWNsXvRNRQX4DFdx6eKIy6gyNyRN3uEC5WRHpUxymb7lHa7g15H23nw
9fiO4CJLm8H2bEbBxfjU0XivSk99SjZtHBFIud6wk6LUJR+eSpKSoMHHTgBkamhp/0d5hwWSU6Os
Lspg9nmBezn2wuZKhqYR7P90nxtgZxwOeHIIqSvApdTL06+pi6/dfHotAU6BCAVJVQltHCl6sBZb
26yi4UNiZ/RunoGw2aCWrXB1pqTDARXCBzk60LcvEumWeV6kjzc+G4UV8Dv+KNAuJ/GCtdDKfmjH
s2HiKC0UMSHlyAi7B2dCq21QUSOhF+Ldo9Tf++bQFsKqrmE2g6SC0XP3+iji+pplR4Y+h9GgpeoA
nAng50k8Dd1FDr00PVbFRN4YyBExbngrLEZYYMJrqvweDFyVzKmoK8E5seS9zPaYWff7RWISVdag
LnsKEutaV66bVxU73c4u5f//AcOg4CKR1xgMd671CFgVIfJ8bf6yisbLCZ4o23OByTu715MQl+9L
JPlXlw/QMM0UXfiuVVv0NjI9biqgwnVYlIW6vLKGAzh1T978kFkeLzukLbtNZrgF8e4RSQvYS4Gd
2OGkEpuH5eU+jr+dG/dzMoh4CPBVM6U77RBppnMoUxXLkWHpkPM1rI1hzTe81yx6mSe2CUUNd7SQ
In2KTiBbOMqFh7HoQRmCCrlAPt2qCeAsc4xI1dbhYpKhZMxJjwuBN2i8wb8N5vmwJHkaNi+T9eaM
xleWHqCDt21jDIxFq3iR+ca/22blfkRvxBAbwqOKcf7086GVRyqCPn8JOxCKLVTVTQ0G7LlZuMq3
sjAZpR+Vhmo9jW3YbefKWYluDgEsrByXYPk/J51WjI00o4f2Ode64rT2hKwfaZXewI/r82+JjEUQ
6mEdpZwlfLqLymKZzlSa2lgNs2WoR8wayeKm6WkJkcTFm9vAa6IS6jE7glxke+i1ubrlneBTq9vm
ajVOY2AMLklb67MfvbaK806zVVBvAr2wI/9vxze+v7L15G4/DoKdr4my5DaMAoXGI97Qjz0zeNRI
7a8JStaxoxCqc8oIiW0FQvK9FwoVLggbTixuWt7M6FBgeK7cG5HNT6zMg55WF+uWV0vD6PToN2ka
R0g00RIVc/f/Jb7nSs1irvO3XpLGDBqCE7RUHvPGX4qNZQGEYHH0Z68j3Xf8Jadh1U2QW6Uugt2i
Bu4lB3zdWIUT514E+Vy01XufmeRGbd5qa+aM//19kq1JArn29EGiXndIme+Fw/XeJ9m1BXvMzAff
SYZ4YQcjbfvLB9iQnvu7JgKQum38dgcXFfpvqt8DFP2b8t/WxU4Hi2GpKfb15RzNVhOqOl/DORl1
3q4r/Y1E4HRmYryuMMiVFPVp+5SmzKao5YLBgrPuHb9QJzxFRxPCOZYemXchTaMIKOfl1mcWAbyJ
/ZdLPu03Qu/hNfkXJrYJmtSZaESMhjxe2dcCKw0/OV54v6MieGfOM+8ShNb82biqCGZdggdXocy4
zLxuxS7rHobjxAZGZ44YGVUGJi86Yc6njQCpTeBJSBqaH/TlY5RJ/gLuXgIQUFriUSqkvXJhFjh1
qwFs3NF/95ELmdZtLBvKXBRCYyeHVjWfsQqkHSO3r93dueSWJ22O+5mQ9EZFQeXKXN/r7GXT/GlM
pAS0V78tkHTqqQJ1oRcou3xfqdXo8UGlwCpm0tSqNax229HXmJEpWfayY+MbjAER2KRfzuNRuesR
+Cm/QxdXcjAEdjMwG1hHjLIiQqRg7P9SEhd079/VsgU2wH6DRO9+MK1skVJYvQf0TKbVOqX+cdxT
LzLTRvzAdLOu5sf8QCUgLnlZRxy26ra0cBxZgQqtIRZotgTzZY0Tn5hDMm7JsM2eh8E8YlxP2ndm
EN4s0qy+Wt6aGctj6laczB6YQpBm8+Cxjc80G57DpZM4GwK2hv1qg0RnPu2QGeju6W//Peen47cc
gChfAukyQgyForKXBt7cZAx0f0lKhI/f0l3f0+aTNPegyQGeXH44l/xOtQsw5mDjqmOgXFXP3vEC
2CSREl+ocrEvt98knEeOC+IGXz8WOAij16dv3gID0hPmZlA28cZo0nHcGMjyeh0ArLurxBy1gG3i
g/T1panaihqSXdfqQO9tDd+PkjiSo16lguze2HoivOhW5Qg6FK04Lyi0PUfAy5F9C8gPbtzjWrcf
xnGUh3ST51F5H7/w98GULOM9rR0ODLtLsAKBgU9X+8nZSUZwTAEYBMEhaOdCldv1FNinWT/7q2kT
88060mpEqwqf0qa5aKOiAI0zwiKd2ie4NnlVR76BK1JBFSUGAPCOLzRhzO+4tLIswtMlY6TXHgMg
znS4xSj+QzMrrx55+u5DkrW0PpZE7pVY4M1PHvcJwDTL3t+7ufyj3eWhoEfNBDgdzCkl7LzNabyr
Z6VLZtnMpSe9GxO5ak6ffoOhs7pXc/4vLFr6CriBzGBugOL66g/hsP4P2lnUlHkIv7rJBFFZ/UbR
/KQJngWCw1aoyvS/K9ioQCSyCJDfZixh5O2quxK+2AgWfKaIRO+OupmEzoHViV6RVaUZz0nTwRAk
6NSddbS9cWRkFxz5ec3vbB8Ig2UA4ONqKk0cVpA8jTaL0UrOLdRu3do7JrVJhTjAh6Bcln6QVeST
VcP00wbAuIoo/yym9ZJkrzaBJA7NTJgliJFqjUcydtzYFCqPUeFIweoZ2qIlffiNnX5cL1pgB/IZ
pGuD8QK2AAA5z+4uB548SNj6NMpMFobLEZd8WH+3WIr8xyezKJksNr7TxsgBdrSp+70PGZl4010h
XTak2EppWifNYB3s7mLZ2DO9BvFbHs5BMhNCxaw+uEnhwrx7IEv4ER6+ZIGX5WeiQiWx5keikUr9
flflfAcSm69S5QB7dK2cd80+ARzD5+jhkOri78RAC7sEsPEXhZVSpm0p541ynluPtC5/g4Bkm3Et
jNQ0iNrB8ceK5O/MVAGZfXJpt/QZNr4aqOWPvKl4PVRRzCRh46ggiDmT7HDulajeKI7LKk8nhGq9
/zsRB2mgV0g7+14AIJkiCh7CasyiW4sY3t4yjT/4xrYb3fKL8780MvpsytLPG5KtYFS3/i5Nwg99
BkFkM2tHEtnZTVC8uRwxkhv6YCxDdXVk2Fh2epAT/HqAreNPTmSYqKu1LQuoZ9PEUVRA8cSh0T5X
oOPjuqqgsMUKR0nACQe/Xy+/UQlawtvXQDWjpywAJdDfoUcmlxXzvn5UctO6wkiTMLzEIf5WYXxm
iOZre5PNJFG5mclmxHvTCwif7vI652a5Mr3LPBn7byLJRqFMKLw9/SkXKtRERtp9NDnsdexmVLPk
UI3+eesgaMR5ax3LltSufWP00rkQwa6hczFZf+LMg2f1fu9gtNCD/dLNUFoM1XhoU1WnuaIUAbUq
s75dCC7Qt3ZDDe4TQmw1bH69CfrDUYeGECZ3xCMO4TIhjMtrw2Znyd5+SWPIRPHzNu61xiXSMY/8
I1OJNsRGQTiCero8g+5eQ7TIrZFM8UGQ0b2QwC3Zmn2yqjW0caSLcfTEUYUTzgRa5rMiaxZmWg6s
TrtExFe5adONEGmWypW05zgGFYSx7dFGSrjmaRRK/Vz3HHI4tMQMILpqhpG8RXCUTBt6B68dLjDi
YLVv1U0dgt0SZgA3qoIk8dKr7dTw1zY0vuxiMTd1kgeX6fh6ALkjeGreVSdPwoJpNeaPo9/Ueypi
EfPYhkXMoXc+sPBr+ozOth95Jn9BbTMSqbW75HqcZTp90J4+H+QMMaXSvs2XrXGN6JhRYU0yFuL/
PhvoWeEZJc/JMSNDVPfwTMNrUWAv1nzkQj4JshvSHkag7QRwbNZpvRASfGyOsxgli6DYl0msutMd
nfLBb4RZKFdEX/sZNanb+MxQPHbVuMxqb21ZSRxW/opaZMIs+PXGP6OmiyVXHSof2h2W4aiDeCqy
B/OBSuc5k4WOJdduKImJtc08bkTi7B8F5JQF0PxfYkrfAmEKcscT2S+yRgNafC2TePDiMNmaO0uL
w9okqVW6zA2703Yd2aBJK0n0qtSBkDaJVWfsPEhB+PDW8NRIGmjfNkB45SiqhS3ApVWp+IoguipZ
c7Lhbw3ialo+87MN+MzHCWy4arD7CtPad3aQOWCxBjVtrvQcx54XN4XBDGxxa+nZL3dKr6iLMI+/
iXFNDULENmpmaR+A3CpTJCeTtD066Wpe/67A5DY3At3qCUVCXGpH2uqZ6aME3NKwvX37G1+4+iSu
vBKHLiIPCQ0zL4zYErKoUinEl3GW6625fRV/hgxVBdyESbdLGqcY7VFebyUodBFFz0Bj+rKdN0rV
slzNTvdu9mfVjT8v7p/1+8CqWGSIA6mER7C2SPGr4A/xN5pW0FieS5ifsu728AgoF6QaJvSDaFiI
CUxsD6TwG8g3CuzS2myfJlnBbRhS1269824kCaB+ZXecz45tGc8P2mJw2QMDPsb0cH2BFkUMb8my
rnac5rlBs2OqKKgJyEGyBpBW8ddXz3We6h+PKuHX4WNVKC5WQloB5BI+29vlYtIaGHypesugsCxv
i/bcIY9HWdMHyzJ+DBRtBpkL3NS2k2c9cjNjdHoamnQ+IQ7zYkiUF1ZQQn2UWuVtctfdmNhm6JUW
rGZOurlZOpQ862d5Bdf/RulGnhD6HrQEzZXHh8/3FdNF+o1t95k0+Ah7Rmi1LP33QKzLzWXsrMDD
/eayaaxm7zmTDSsbkOXP13rxHZQGWrqTiG7AZwUCiVuComxa/y1lwya/y0qugIo3BnFjVln7zsuo
KfAlHxqOk+SpAM46jAw86nqdh58nW1/9keAKiPg6QLgEwhFwgVu+OKSXM06HJuJFHDBG1bX92XRF
L48U0Broq/h+JatSB6yiKzZn5Sbb5p6RW/9+EFaOLZAScT7tTGSXu76HtN6/tcYO+o5H329Qt3s9
fMQvmTDCWkDOFi54qi8QnRzJKBns0t22e8X7YrnPNLQCa7iDg5X9xSJnrSgDJIUCc05o/+lSLk8u
2FrssAqz3QL65X8IJeXxD2+xclfUqMvUUgkyzHjBfi8eZ8ygYreClm4t5IIpw5ibbp9bO/SfDQn+
/hN1/zsv/qKc3meiK15G3ycCq9QTfEW1ePhCOQFkSjp9yVVpFiCnSwCXN6Kq/j+kM5gRn5EzPxuU
qCEAnoucBb5Me0Y9eAfpsgqX5fGCVLvM/Ha2QZ+6b7KNk3NAO8FEKtv4sXBrPoPaagD09zpOhXRH
q4XCPtU53lgp6Vc5Q+VECGGdRlA4zA6bosg7KM3D9y+evk5CfpfPznTMHpxVHD++4REm0sfqxkED
FsP1aAYkL0dUnh9wYKiwVEgy+ihw0ID+MzbDMkIiHSixsIZfr9zd8dILjK4My82IzzfnH7FoU8Om
+91S0wqhe79EnbJajyKfanLZrpjNCDmL0OXLOsLMFerAChAJJLkWOl60Zbcx5GkavFSYPzwzEkuH
DrVCAyXrNgrF5dJQE5m9gkCRkFTuLcjzDG0+Jh1w2HOuqKYU1/L3+3W5fQFt5Qxa18qO4deHvwCe
1R4KusYfppibp23/p1prP0T67kKkTdakqghHOmrQQYM7MbgqD5RSLBgn7QC/cjvhgUi03CLDkCTI
aYfCExVQWdiXQf47OFccIObn2IEMoH/d32xHBbkP/Np037hagLYsDYVY4eJqbSiQGkNV4hglKsEY
w4QgEcfvTiKRtW113kJ+BSu4UGRI48oYFw3k92S3dlOJ30wesHxyVfpRfi6jV7i/3HylF4ZyHxCO
DCiaNoxqYXW0mH9W8ICoGetpjSEZJfYiZEhGs3A2omILMI9lsglDlMv/GJAil9wmRTT3PuieYFIO
wcoo5HJVoK5rJgRWVdKflf+qNp2iyqOiDNNvDN4ea2JPcDZx8dAQZQjatDENIBjz/meDKIRpn5BO
5NGZb9fHUUnlWriRxCVXEV1t+0WzlvYmjJXxPRhJUXQvglZQcXZ8R8z5D0J7cEfaaRt6YwijEYVI
Suc8bgI6AijI4skq8jNUCDVdgHzMVj1MqrOTWMKyMpZK411svzV+YJ15ODAXnxCsKtnV5NehvT26
ahrxBSglHC7Z0kJPBcusEXbE8v7dGrw6XwcrytSe/7MouOj0/E3R3XqiRoNxH0lPKP5GDKqq5WBD
qFoRngnQjOPrHxdGERuP7JiQwGvdeEQ/UIWD7tD7T2RMQXme7x+j1ovjWLAFybZR2dT+hAkr0TNa
cWLxJh9qIhN+QhIIwg8p7ApbB3GU9doMLh9MGjtCPUu7uXalsL+K73Kr0lGqeVYYDcdZnLlBl7jF
VzEYjavhXn0itbxmDqEaPxyIwDqmVsojkVgkNHNd6wa9tGh/ggXyfhOdakFGeWNA289vrnHucd2f
Fxo0B3BG1E7zt6c2iC3EYlJfTFF/D5EOmuXTX9/h3jYqrfBad1NyY6StqpQooynbhS2Zc5OpfPKv
5+wTB/NI20jHeNBBrTWbmQLx1hKbPCy6Eep8Co069SOqAFcRY+ocbbey+kvT7bqV8sqWWJEv7BpZ
kHOhvty5QDkYOdsuV4iFkX5vGmX0KnjjiISmWK3Mxtjdxd0kWigxn59qy0PiMdqDRM/ZJ4H0Vf5i
3fEFYber1vHj+PsNBS9oo6vLrSTKCLleohlm9kCJbdglaBAHSPCVSQCow+a9KfRnlLqZcvhq2atL
emLaHi2kROsJWj2eUnAnW/qD2qbj1Zu0a7CczaVKQRvYuZecVYKdDhwL5quP7xapYPJF0L4r3OBc
8EKj4TQf68sFyvRVWhnRJkL7AmYAK8bog02DD+xBCueZ7eXPcj0Asph4PBmTW0jmWpeOVZWgXnzZ
77ujaIFV14VVLWk0CYr6efCzPTJOTSPYVdKRC6GZ6rVXoNXrKQ11/vw8FYPPNQDTO/NJLhYhx6tN
sEWJbfYN5hta0YYYTluy6qirj1C3Rw8El6+UDsT7UYVOu75CWxeVN55It/k4n/dfW2D9V3vde8DF
nAnEReJhYlo0GIWW2xw3ABh1CwBfQO64cqirlop8vIADZW4krnXuYgdi/HBKI9qusK8PYHmFX4bu
N30q9H/6LQdfI0FB/2y79skJ0vko2AH6BgM+DorBul3EiTytcsM47tqzbWA9OC0hJBroGHbrXtGw
nYDiXRqM2JHYAFAYWZFXbJBDiQgntI+erDbOnvKvX69DSlOyn+DeoxDMLqZXqFuVG/Wqd++plZ9z
ilaWeTH2LI+YhoPPtniyyd25q6eSw1AclRFQXNUNBpKYzLRHkjr+3zBWkoex1ZKZv0GBIZMC5sk0
V/tJkgFEmDy6LMiI6rwHCAP7rVYfbdQUzzAiTfBmFxEfisBsYHXQaLA4F0nHsUKguODHUOBFvNFm
9YhAjmRmVx9+0rpdyZSGvKJpoJq5MIcScrVRAW/zfOndE9YKvTbWkwh4O2GTHgsUukXax3uWrmP6
IruVFG2cclf2bSBIA05JF/DSA0RJUazQ9d+voqXIcCHbTz+BEoON1r9A0o/L/yPO+I7tb3rNVPIQ
A+eFubYfSo15hFTtTARjJIyVkBZ3OlF15WnmWLpJouoIDBhPRJ9QfQ6mdwuax9R38pZhLFiWShCL
SSWz9CLEMzwgc8ckyBboeljjWFmSea11PclL9cMuLUp4AL3A9c9oHcxq6ZTPcrYEfUd2h3okmhnT
YmGmC0m9QOO+CZKjRtcZZha/mQ6zpHehLWcflyQ4Xj+y1OHFVOM4MiPoNWlP7SShWPRItC6hWCbH
biqP01qpURyJaDNTcUfD8nnIa1PaDF+JPDTxZPgJ23HbZngTEnG8O9BYnM1JYWOos+PpV/85r4F5
CYmTNQ3xEozvsK4dg2I1ANTUSp7mtcU4qfHorHjSEuJebwu6n2vU786sLyRoKgHM4fQCr4wRUmvB
4JbCOfanJScYTCAJfwFAlUvIEeOqJaVQpZxd/YLVIZ+IEtteFJteumRrG+NYPWB0+vqDO6gNvB7Q
QoxymH+JlNAXkgUkE4QeZhliTweVj2RDUtrY5qP4sV5SHmRY5+n0vJAO/gIv8GJrMhp0wRfSxbci
Kw4RFPiwB9TnbCtAGT5yFuBaSB1vtf2aNgH0EgChREpYYf+rcern99gK9gYmlV0nmi7Dcf1HfT6s
rUz4D9fQP4VtRFFkGWXcC8VkySfCqHis613D3IC4EavaTulNOjKoqSN1Osduh0txW+uQt23bKqA5
Zwo7WinfHsvbAGh/2NnyJKliD5q9wlvFnwiyCKa2u0+cStIjO/in14mDcLncUfn3Cy+mH4YW9+gw
VKfmyw4FO0e023niJ5bxNMfsMwLMZGtobmkHNWj26WUeZvsFnRNLm4Lao14AZDnYsfLxmFBHpAmI
v9+s6RUgXebDrDVSqalQe7gbdDXQLjqvi9eLtM66kz+rypkTRID9Mfj6gpS2aVWUCPJG+7A7r25J
qCxpeEN2wzrgsBC3UAiCP2vjejqE+US1oDIcFKsH7TocSB4a4hfch6sH8oFmXjVUaO6eMVQMlHtO
8QBEruwEyhInqssZ9ZCEhEjsQNCg1XXHYK9RbQHsniHEGaGzKuUw4Z7/do4gIug86wpb/0HpoWOO
1VNKutZTXis4kAqCa7cadCsmQ1C2dV7YFHM89a70vgt+E+LFRliLIa/GUNGuD9Yr+a+qU4e1nmcB
P7MruMsSYw6LVLMhr3fC9kvbKYHOmupc0ypxBFJqIS87QDI5PqOLaYgisHEFtFEQw7n/dXkpX8j1
r0lqczLU0SarZ5dKsyXAYyjzzHFiN1lyn1gWdCCZBXk8GtkKMp3yHYT5iIroHu7Ro8VYtFI9mNQ4
KLRj4wqEKkuftDH4tAjaUKyg+6DsTemZUieEcAzU7Pb0ylOujguzwGJVbRgAk/zK5YYnvtYXWGj/
INsRhh6PmJ9z1NRZ+WIDx36+voPVptZdhORHB7lQh+iSeusUtOvnBqLjLGnux6gRrmr/4TYLwWnG
dHFYjM+oF8kFGeZyxSIj8gjBSsmuHY4C5/huuMonr/JwZbiGSQNhAHELqGNURkLpUZUrJNK/UzLD
CLmIcG7yvrQ86S0MfXp3Ny6cAg8Y0q3sFXclRAc4hwBYCEoQn9xkJJqIHEO7HOD2fvvTj7PnK045
HwSECBzgieryboFjSxuROpM1f02Q2RU+PHISlfrTp5tsXk0F3RC01U1MxGK3qXXKv8mzeKPxDa18
4hmUE3kI3njphaIQohLpT8Rb8Mfqmn0GGQw9bc22dBzViL1PD1ZqUQWKWaE7Vz4WSA1j4vn82MyC
raRiknUNH1ipP5GRpM3hkFC01PgT6W2fwqz8LlTy1OvIXT14WJ1VVKO9u3IDk9XO8v0GEgvgHJsT
kdMrvbnujzxjLMBYk1ZpxSz35mFWMASYBGJ/lPkPMFiZmM6LMMZQft84W+E+I5I3LtWHiSox4HEX
SFuG4Qie20VsEguGRmx6CJd+wLGN8j5t8MKHg9BTJcV7BwFTT39XrQZSCjO35GMb4NugRHPD7F0m
mj8Jo4EOFpOU4swcBkqvtQqATI73HzzPX2p7fwtwBRG4WlGi2v0V/0vHoxPrnkEMweag/YiEFEga
F5o6F+O51Hwqu9KC+n3KeTE95n0dVMW5Db82qU+/2hNA+DsXEDsnWXkLDj9f/sxgI/J6Hs3m7+fi
AeS0VzRNZkNjHcZo5TYkvTSeGlQ/9Nf2DM795itzcHbRtQKmlv8Fp3JjAiRJKYBtN1J+bvQvKEo2
+0frezIqkreJRSXO5BLA+fyKlGv28f7Ru0jkfzj24yx47okV2FVCTMvnMjzU0Mwuxo5/rZnDTfu/
gwCUHDEfFdyiO4ut9SQmibWhXhXDgPqJAzvECFbbwPGDnTfvYVh/4wj9dwa6iEWwbKfseEN4wvn5
VfNsGF7yHNBCcnlUiF/N7p9Ao1rLrMO3e5Gv/NpLApczIsWsP+ODTTZZzWiu+Kv3vxIwF+zUyzNK
oHSiDbnxiASEfs8f44DBHJr9TY8cnqAHjHymP/BTYO1Yx5rORORssIGL7cl9IojZsSzuMt/3OuZ1
pQxwhMvAs3EutjU8CNRyLL5FnujufjFcGk1fSBEJGw/9AhsZf/3KR7/uykF9Uv1Uf2b0Uo9GR/K4
IW/UP74H4emNoo0yZ6cvXzUkb7CG5AGXz4aOtmdv0vhAcyNpnTZiXHSgtt5ndp/3V9mpG62UwPpJ
T4JrpqDVy8V+JJ1Z6D1dvaZup3P+Z99wcC8j6cppMed0MXR00nyKCxUgqXZ2q6FGb5BCtXbYhsPD
LCZG+NacY6fuoa4YCi1eGdt6PN7QTqD1qNElshtMcf6sDvOYrqMV+MiHyWw7HHJBW0ASCsEZHPfG
GHDdnUtJzsUSMn0lwvFclpocbgp8xfQmtI4knNNTnEWzOTcm9rjvjEWjFpE7hQAdPnwS3h73+W/i
6ijs3oJ5/Rl+wEosrfirXvzKlVLiUMARrrPjAqBccg0flLNa6pCSKnl0hXgWlgVk2sgnsLvTploj
fk9wCEJT9EF4Uebx0KrGo+5daE2RzVinSi2F4kRqzPCtw7YRBI5tZ7LkyU9FkZUY05/CS7zZr9Z6
jyZxPqGNvSApUFUUkhyqlVEk8XejABomhq7AulJIOG/2/eF0sKc1EEwfoe9+jRaSNuXZTWIxGTnk
FIn/eAqWXM0DaZNOcLXmPsDWKkgHepSSeUJHJGOGcmWS06dlucqWlgFi9dP7d/17l0V/8c3JJsdf
jEGU+EThoPf/z9ARxuvvKJ7OQDqWOr9GfAZOD3DJPG6aYdVvvP+egnt/rSEcWFZENXIt5B4nMwbl
RM1afrWPdhsiShkpUNp34erY/4tu4d8LBEs/GrF/NkqXv6wEbUK68RTz3iKQuW08+RY8A8fppF/b
avAK9QtdDqILGOql51zqg4emfxxGjIdf6O204IQGmsWABmA47dVdnCGDeyoix81Ico6u/Rlikayn
MRPLRH/Mfermibeh6dfTQkCRe5/sDy+HworbeyUwsZhrX0XJdGGzUVidb52NlmH08OnAGjOqdg4z
DucouIUcrLRd97O+9wuFpTWgv1Kf8KGz+TUt2nNGjxKEKe/4MBDceBTaGQxEQIGX3pvel589Eh/t
VjIeaBAs2CmUt4t15kj67BcpexgQVV8a/da05vpqIPLQPzN2fVxsTpvy5LIIVL+4lXGtVRCbnMWs
P0oO2uH19DPFv1eAe8i43EiUcf2/G7BFDciNOu+R0a1WWRWldm8rvCSq/havFTs0viEH7i3Aw95j
p3C64FUmcMw584/JYk1A0GIa/JsmWzT4IPhVn/g9Y2SetCNnvtG7cwdJRO3eNMJtGza22kixQHuI
h2QlDLzxUHpSvKOZxcvFMt4XUmZj/E4rKfPBbAQTLNhG4DfVcEzlVjcRmcNULKdw1q28LbxaOhZT
fEnLZI03puIZDKzLFy8gUBCVoGz4S7ST4bWFiV5uwvGvzdP3vv+xy8hTFBfZ/OFBHfp8MlkVpHW6
QOvo4qAvcC7HGkoEyF8lbPKoAKzLR3KB7svPN3eEFxU8L91hcBWahdttdODkYZWJbE65uCpWbDW/
iQC9fqT5qT0x3t+i1MJ60xtbxpjbN2Cc79eD3TAYnEPJAdpiWUUsXl8EGtFXhuly/JKdNsb8i/AJ
ut4MD4d5PdcF7D1Tsa5JnBNW+Rjk8KkTsHH9cT4iHkoP7A5XWCbK1d5vJae3GOVba70tyXGdMCZy
WOx1oaayR76WDdX74rZzdiacLcDuH04tng2m83A3CZXZ0Bf1UcI6nkqU8zqH8tDzarMYIq6HZvl9
qIxi4uad0nNG/XS+1Jo4sU4Cq7OLFtithJzHMk4HErJCFGp3kOD70iO8eLwl3L1Syxvnu0AKs/GP
6L2c2EDcRQQEz8lWwBeco9zRtyZcd1KhULBPXdz0V/ucZsJCIssCJBmFua8gOYO2z02esVinF96L
WdZcbVUL5qfnYE4WJKGQJrJwutNFnLDOMxqmq85D90/XubqS+TYKpLiSL7AVYm8UIYBGH/e/FLeY
iYl28wPG7etYxA/5XiAf8NqcKBSGjvF4Swevvvlh00xN04JHGGhhnYQX0eIj4pSHNIsBCDBDqVvj
SRNWFd1i9pgqPzdw2cg6AqoEuofb+1fOS/l1ZwtnHwKSbnRkQZEOac8SkHf5lXCLQISV5tcJQzcc
PDLUXRZkoSy8p4QrW1mWnBYqV82HL6UOUtm0AkX4MS8aa3GY+2B2Ha1GIbrfDuipl1gdGbllGLVH
8IDt3uV++UHuL0wWUzRjeW2uopfkxlPEooV5yDZe9fzD/mzZiF7oVItx6uWvWqPJmhMRG7qIM9O5
eTSqTVX/DK2c/sk0H8ufa5ZkB4iwg/z4E8gZQyBjaQJwaYbiyonXwnGKSp429BG4/t28bXEm1QFw
iLPmrzujnNWe0g7qn28fc+DnwGU1hKH6uEyFUnzn+U4Rhsyu7L4ERRD4mzPjwrzPPTvMnUr8eYc5
Wv5Ig3jt5RXgtT2mbZD2NtQRXdJ4n0hp2bNLfhlsyMM5oUOB0FIWSFWGqfkbjLBPpE5vnSM0TX2s
7NRnLuNTLyOdkIW7p8DpSmKsHx7NVR8u5u4Oeg6Uz4ZtpvI1YZIj5gT8rjs/EGRqTY3ad/vwl09F
LDxr9NjJIM7pcjFDDdu3+ee5kyRG4veQl4PFcn5XNkCfimQu4MUEvkXGyCgEekUJWFjem22LJMMN
v5VQFZPEbjXTLTSYuGa5S5ZhAAHmh8C82iuHjb1UlGeXispmFJ6OomRHTMRJxJoH02DAkJMxEkqD
S2SCMVFjQ20F64Zm3Vo25rf4Nl64iGDlm2dPcZxWOn5yM8as1XUlg8FBlq8N9FyUDqelHPAayUGi
x06+soTiloxZ6UTYaVwpLwzSD05hhGOk4cjX8O9dnfknJzMUQXJVqUyInH30LnbHdOyJGdwxh83d
6bZgknQWHobZrn5irYxVo2kG1FU+i+Nr/WdbMxK4EPlA/MwzvUkFwiDpxXxvggvEGxT0iMSyJ4pL
o9OiDt5bAvcPhzQHZ+zTGNzpCtt4ie+u1XU1TWtgsivp2GF8e3N6Tq9k1x9QnC73HBIudifJBdX7
XXX1j+Exwr8Sadfjkzov1Z1oLQzGJAsRUm1g9oK2FSRKX+2xK2u11GgivWwmfuztQ8qVr/OtSjQ7
vhzwMRgtZn2nPeStQnxHvH331ByrFTu6QDupEqgkZCOFrUEKpVhwLVd440AbVJyQ8/gjib6JwdOx
IySYbPBpl+M3LgrOnRg7oplHCzdVXTvbE+qzdnJTbat4shHtXlMyNbZX361+CEGE0KCFS4JUgSQ6
VA1AB4bPz0/FVKWtOdEC71LAVVe6G9MIQZKOK9wO6Alg3/R0vu3e/SZDIqCP6TRy+zyole28bk43
/GJQIPP3XFmiUn6wuRCFGLmOPajtkpqQ7Tdz7oJiC9lbHcTwAyDjmSKjkkjAr5jfIKOT9/A7cAhg
u+T0qrOBio7W0RppAdWvKbx2RCCiEu/OtPZKoa3IN/mcA08PALbLnoH0fPeF2+Yzlqbm1OZ28gRo
JMhLTgPO4lpCkrGnWhHFwptEWxxTB8nxAGicLL/R+/MjE+kMIXOwMUGQUQ9+GvYnLjFQ87EYVLnp
k08SZ4KB/Is+U0tVnVTfnztM9QfoKBcKlUSbZCapzTIj9MXoE1Ncl27eN0WbnZqM3R4EK0Ace+x2
h5gQ6kk8VP4a/IDxUCX7k5KCL/w814bI4bcDLjQ8gkBbRG2yLfUz00b/Nrb3b4llbh5n9TtbYnpF
olwaPCuOfCmQ1cVOBlyAz3b14SsGrsWjPbFBmgNtf7oV1042d5XayE47V5sar2BsZbpMtclYoUIz
3EwksktxjrD6bzqrQ1wsRsv9Iiu+JqL+yGNHfGRnBRG3/w/RxGs/4m8jjkd6MISIIucssR+2BM8Z
CSq3531YsHELMZEdfRHzxpxamnTDXn4wOBbk41pfRWwOJScwLCI7DK6YeSCvQKPkuO80gFCs3owu
pI82K7VQIsZWWOVqHc8/W9FVzCuz2SNb5TQDgIUDUXEQu/2LCacljq31k5Cqcmbia0AwA7L2WDUc
3ymokwCxs20YxVD7RacTbPqdd8WkzHDbB8Hv6ivAnxOyYgL4sDnGFUmt57XRW3cB9kZDEVKOZg3Y
ypf8Gpgk2g6POQOzkGw7Kz3ZWsK1zcPUyDgA06eoywp4qguAn3jQyhrQyAJlBYSnwzCWcaOf74YZ
kKW3SOiB7Xvn9CuAq/X7i/ICjZsoMUBnYCbji3cuPNN2ElMmbozPUoLEJvd9QXFgHc2YHP3h1MpF
JSpRaKAuyeKkDHOVwkuwrUUqJSghmT5owJk0SNqW9+u2tElAkp+mObLmU8kB93pZIHzadzAZylVV
mNNaHT1V/6Vsa8g31UNVH6dsJVDuPxiYdN+LvUQaQDM/hlvf80uZAhVDrimaO2N1h2CXzn7EnsCg
e2gj/fuqBQ4KS9oJZwZoDNvG3YPt0EOTU6/MB7lK7+Frt8Vkyk1eRc0NrMEBkGr9m3dscJ/JS9Nk
PZ3JY0gtijKszAsj7XAlCp+xD5mO9hJze1enNIHFx0+fmlFI8MGJNmDKIVe2XvuBfEKpicT7rUhg
sDwyGaJQxmKr2Q0c3W79l4NGCOBuNnM1K4G2M6rGp/z8fXcU7I/nNuKCLN168xDqfg1tvYgNC9kr
PeOLM62UHuqd0ECTaigwWLY+GpuhmruY91Y/kYAOblY62/7MBAYlncKefwUoazYEzb5gK0GV3BeK
NYp91KyRBD43fHmDWLgCzyUmYR5NyRoj6akSNx+mu69VIskjgsxUGC2UjWoY4iXnETSqxpfZ+7Bt
//FQrfXv/V/P3g2B5f9hAxecdjW/vvqFH6rv9Ks2UEI9f1Qkc/OeWx03G6mV1JZaZ0lVD8qMGpEv
3Ep/yTTTETwARXHtzGwkZntGfeZLpBl1lTkEuZjJsIJEXISaqAzpGxVekcyShWSMC5wNlbcB0MAy
HsyXKU75Y6rbypEgjU0nR3Q7ei10xbHB7RsEBCAOOg29KnO7s4594laqgfrpjt/HNcOQ6fxPh1Fj
N2uMvzlzhjbyhDm+FNIlAyOlbUnJOXeEG+IpJUHY1NcL+bkz9oEYchvl70vMW++qaTpcDLOkc8Sk
qNtyZzYysVp4pVJuMnV31gm4LA9GjJc94/Y0jGLQS6G2IRmOxY3SyysFTeMecbKBRL7IUrfRnUMY
o5swmceA/3/gyCoeugIly7wSTWEgfW5KBO5mZlD7LloCdp5rOpo8qhl8VkA2Sr+7MbwtsBUP7DIY
qDMLXTJ0bgECQP+TDEX1JbzNMT/pB8q7j+XDxdETSt9vjFC1HDFRsSqikFD6g/gZMMIsoAeAf+u0
rIXkeNowNSdGZRAXEALGufg5CeXKA2/Ly53hvlK5UxDJ/DYVs/M77Bw8ZNt4Fc2SYPwazBGe1Pmj
rMcokhesqNfkAxNQ7xvNj98cgcVFvu18v2TUozmeCcuz6adaZ4FUvKYzwQNnwUmEuo7HJbNqLeTI
+4+A5W39MQ9YX81CFO8xflXQ49Sa1MHQwBJK7osZytBOWyjceTYglC5ZP06XoLyI0S5qmAutHNpk
s9/B7YAu9oRqWu50e2NFX8TCp8iUil9nQwZhkKebcAIwoc26stKOHAm0Oct6oNjx6L1Whemv2pjq
CNuSlIUDFmljTeBoKx5mJw+WsaNUbSMXgJz8ZkG9LTTlgajLqtp9LLZq1WpJiN7wLTy+KjcYvacl
mbtjljdn+vlShVDsJbIzJjeSalnFor4Nt2RZy1aAL6BkrcViq7WYzkv8woCBGem0NCRaU3+I8f8E
6nIExtiaj1bFSNiX0uXsci5kW9nmrsXoP5SNSOifrPUFti3wuVVcafK+zNjdWcurTY/7syCMrVzI
FWoG0eIem7GSuQ2VPXHabUTQhlSExkQYd0KTUCsyDjQy4Mq7l+AcjZ5xh+1wrM7sUcRiWunOGnIX
fZaLOw8viso+pLOYSrN7cWv8CVZ48jmwD2RVOIV8eCjpCFXKaIn0wl3KKZl4kx177HYz4YNNTlaU
KYEYyLPfU86tXAlZCo1iXe4obQCj4UaEF67uiAdVKspMo88ZI7Ks//g7ZXI0l/uMyGNNiipIZR+F
Sqj2Ql86zmzsqhUrLwODH29lKBico1TCozuN6s2YNTp12AzHjzdI05wt8efVC0nEGSOLgOgYQjoG
k84puH5O0YN9NlGv05LAqaus2i+IzQnuDeNX0Eb6fj8Oh8ibKJFFRWKhwsMJG0/AdVvPv4LNe9ep
0kclL23ZhfX1Szx1HJv08RepZkmMUGVr6by0smg7Lz3+gG8kIXWbAH6IRAqz/JOHgJAKHJXLSZlb
FKhaSkZLPCSrXtyCzfGsn27cCn9ZXsTTm3ghATrYZrvZtywGU5L2acq205wHD3xYPAqTlf2DVbh0
e77xb2UIrsucH4FcV+N67PidQdoIEcAPfRN+kcfdy4nL8Fmc1aHjy8W+pCyBHfPlp/vo2JpBEBJL
pVjH2Y1WdiEIv+38omxFmhjn97dqd1WO8+oitfVk03dki7/9iYgHDo/CWAOVDp0z/xkBqJzmw6JG
9avoHzbgOIACUXVVbFQKwC0UChVBUl8u2+q/z0V44AhHvz530QBI5yjIMxe0hZkhg+lQcZv0ae0e
eQ33qgOcPHJvVx9G2b75DRiAlFzUYe5pRb1yvHSf+MedN6AnsNigGk+EzVTrEWBnD/eHN4Asij/P
etQwn4ZpfnMvRBfpVp7V44exEXBjDRQYzWR9jwa5r0y17i/oC5FKTjI205r8TDtV5T5kg1pPrTTF
m+RiBmOxqGUNYIJx6bppL2LqhCRL9+C+C6u4++QhhzurMDtNFzqpWQYwgFN8uPRgaOET0N9rnbqV
FU9fY/DXcwu9BJuntbfYN+LDFC5+k5qEbZw6AuVs6LJosgtmP6XKRaXTIwKaOTMbrv0jv5CWYL6K
rw0I/oUXsiFMwFKPNwrUZsqJvtQG7bYij/rrxlPDj0+ppZNKRjc7TdfMa9j/vPpx7+RrXmK6zmiy
pEDWISbNYOP4eiYhs1rn3hGlvWmASRanUfiXU19rjHtbeL2/w+gtDvAT4JSUQo1ffNd9ZzU6YwgA
sndOBc8lUMA5S9DEpF0pcWJCzRuZK6rrwKseNZ0oq8plmaL21Rfb0BIv3J+mp102F/8GlfMpMKYF
Ns6pOK0RjtyWX3Ci8uBZdXZQo1D96iOJffuy6PofX5BJ2P4gA2Ez7kvKa++Ih0GgLzGwIi5K8PFF
QJLifsBvLZwKfRESosAzp2uX/pLL2+gp/EQu6mr7zbLKLAcIo+XDNoI6gT+VWu5nrdOtBwOLOA7s
JaD4J1o5W7nDcgtRvkkgJMLUCPi++INW9ZeHMBo4mL1+mZIDjZhA7dB3g5PEpT+rqioMRaKacAkJ
U8226ZrNoigCQl9aw8gbYAsGca0E7F+MdtQJS+k1WDs4ZvWXz368yECNccLjgW+bh5FJoaJOCmWw
YwdPFrT8nU2IGMalkU7W/4T47o+6P4SOwsbxZkNcdPb+QvBYPeCHDY7VPEFnat1DhVz2iUgIkFTO
Ly0HYZGPvF12ITv9fI8avG59Wfg4+q9BcvZfrmhQ+BG7+iOALiXNW+1qXoEMKgVGDJi2/OCI5acP
8eQTE82G8RHxbf9OQhBfTyb+YzEKPjLHVFFB3L0DeuzwHHIne7XBQtqjZgotjzV1kvpjLG0qTl+r
51ktgGILaorwtbhyJG5Q19Mx4zzmYG4dVVWWdVUDRj/MN+VAUrmBkHpGcO3oxPQNLT5WPeTQJqq3
DOECLufRziESsuwt4lN0q2y+8NR7+/QnKYB03igfKP0dzpkkEOEdmzJCiQj3chufdFqvET4oPI5w
RpzAQFx+Od1v0tBQ72hWml8SRwiTEPW3rwMWVWFJ3OfFo10YM2lQtpZkzVq/RPU+09kJuafyGcJi
Cr8n705NkSO1l6LDvIcYGwuH/Mrr9mhqEEsjQR2OkVNdXX4GLK0xcJkjEA+Jhg7yRzQ3tnbk+13k
uBT8yro//bSy8mw5Hs/YW96VusvEhZahX4+oq60kQ4TrYgmGAmtGpTR70IHdcWtoyd6oCJ+UP89Q
z9Y4WANF7SVzpRgt+ZjFjnm3Nd0N9u8daKH7hsCd9Ta0X4nSg60wscv7PmmvYnXILaNOVQC1zl4/
Aruu8fP1IR/hr513+H86WEg4LwAMxkWIsq50lUhxpnSoFbYC38KWs1gHSeZ1yn5pV9ee4KKzxe7R
1s/3pkeddmpbioiflwC/wmntQErYqmctl7ON2zx1uepY/3jFg2+4lp+iNK2kx1sjpqt68H31p5FS
ptELesowXyumPH6ZZOaC6tnvkALzkf0wFFjQs4SdMBeJTqacE3lSGFw9aVcTOoWCR5iG/H619FLj
qOByaQvREeXLNAhOj6mSjkvvZuW9oN78bZ8o7pJ/1MH1V2xvuBY8BfRqmszCLKBXxmy1HcqG32pX
kQl/jAvwqQ2UhBAZv0hnz+NcKiU+KIc9XNFnTKom+zrde+gyj7SF+YTNejgM6X/BiDof2BKPi1Dp
myPWikUDBJfkQVf3t1qQEtdC4fWBVOmPBMxUOjvo5mkIjjeXod24la0ApdDRvp9IfYpN2+pIAFa5
4M/hQ5SG8sdc52qaI+T9xK7mxjB7swjjTtgLhXmiDmh4HNptBxPgdjqZW/VE/YoQ2FdW+Ts985Nb
+ET9i/D8LJHKCYRapBahRr1ZDBmICufLF5B0EbPxnwuMEoAYwvr/zNjcDKjozCqMtA8VtUGf1mtj
2rIcOOGMsJIbfnvx2eRECc8/XiNAxd4bh6IGQELpa/2nPCSZHF9tuU2Bbrg7Ub2fRF7HvKzHy+DY
gYFvyUa7/Bzd7SfZET4hYcLaqMeeOl3HWL5a3QBqJchw3SP0vWx7c78PQUxBDldhzOdrCYmghc4m
qjqI/TLHRSU6cMvLGAHpnhWRaQID75zkN1NfFamZr+IZpRMFtX3KhlgK8OX4lp9VDKVl+1Krh3v4
gk7u1pRkZVGUHnGKF8VaJd5LJIyDaj1Sm1lBl8DGqCSM9vuDEB/g+pZU8mxhS7pGFr2GdAuEW+k3
ljtKhVG9urNMYMziKY5ucKIs6FpWLZJzW4sr1wRP/AXsyDLMqTFLSxI2hr6fz4r0SNyfVtCCD2p1
K+iE4SREGElz83hWoUftpn7X8PQdzRwddynkp2krug2QrV8qNjB2N7bkUzcwY9QKfXLBey2qM73C
P0KIQ3WknIR+v/kkMHP2KjLoOJreVKXExTJLka9TQ7aj5+nubVlW2MaQd0WUSBUbZBKYZC85C38G
awkvgwAn701ccKMXv77Acx8bnYwoG+zIABg0VTzBKQzBcfkCPXQp4Kn6LkmKe+ZPQ2GhyRKDWRes
7GSpGXhldyFrnNpeY68enWx9UwxdKMjPtXcOCgq/deo/xm7U6jEc7mZ9X6JDfHx7pgJTz7jmA2s6
qIMedXqvmQXEDeWrPXvquf4RJipD+secRAB6eqhWUQI000i+bPgy5HCgnR5xqI8r2ggKdmMd2dqj
wMA+H67LAxk+kVT2Bl8cyLyEE4PPwKGjngZzldi40ikxVJ+72RPpbA8d9z60sxGYcW3mU4q9GX0o
7dosJhefTnVIadhnamYLAqw3B/N2R+lfpO6sKJZYVV+eIWrX2vPFXo0z5HRqjD6T1DU4MriwPH+M
fT9YTqQe7Qn118rVhrYQuoIcU6nrD4JT69vBhwibsR/DOANIKJ7ONtpKGMZliiqYMzt1+Yqm5efi
guUAm1a8nr8Shs/PL2HEqpZREO8WYCmOjClxe7viQHYMINofpmzxCaRzTdoJIEYXFuR/8Am1lcpX
IHA7swUJsZpCQIK8VFQ4vZOnR0u2zzxQC2fRC3YY+ZcGiNWa1YV5iJGYlpgc/0arMN4msAITWnF0
qqqZitmUvF78FWFrDltqsnbKdNKhL8zcOrk7pmpfUe8FNG+EJ9AN2WD++dVMlVfRda7NBV0BNB/7
pRMCVXF63yCYfHTo8iHB5LlUG6eFAUQROG0qf6Q3bUkUJBLXWKSp1nerMFiyWkQ6I3hTU4x/exd2
Y2fBL/WPaEB9990Jf6H20Mc15S4xpDOmOcwqPMKWlShZFS6FqSiz7Gd6xlOVfZ3xgscb3m1jJ8mV
i6oPG2Otp3pJapS5LegFjq7nuEyPfk9jeQ3NmzF2SMiE942P3v7W9b5Dv7ijHBnCDshU8ZcYkNvf
zdtAhXkU8IiimQqr6r09gpHtzKOvF7WtF2QYom2s5MjDojyA5HOR/Vh14cKE4tzKqa2EOtuWuqS2
51blDtOEP1BE38t6zEQvQAu7tvHrAhu6Ck6cmmIDwjTS6FzJX3S/L8Sud33cQdyrGE+A5HgtMxaQ
assQhU7rZFtM3K4CXrtLIS4ELC+yztdiTGSdNXXs/InAwwPb5Q7k78YVNnugE1vkJhAtrr65pZ2J
Co/+cz+y1ue5mkgXwGQ9G6McrsF/RJlGkiIUmYSRcATu03uUH+rxWV3zjDTVWFvwuhxaXR14bAWF
amO2qfudu1KvtWjwOeJhI/CXXQPpgzQOocmEyR6LPEonpTdlIEfWFSXLYe3x7GlhOiszFBf+xgTr
M+erVifZZZ/IkigN4SA5g/x6xuMCaoE52Ng55i7ivku56qxqWpcSPO23yYJ+MoDIkWl0cMkmxIQZ
0tYB7ugbrn5GiMaGH3pzhDOqdZIBzHiH/9xkwmkRS6ncEMzPwX8saPNf+FK2Ycci++2TRAKM6jSD
WQh7MPKDZ2Lst0HCZwoGGxOpgdk1hZyOJi4H6oGt65SA2eoF5trvJVhs4NOhsU27vSWmlHeRtece
iFPv2Qk0Zbo1P8yD4dtsOSuVF8bt/qQ37qn/3FYxaVJPK9Qsxs093Z0FOPnKczdP4cfA/4DEjdre
PdttgWsmumlMgTzstCRox18wag+jvzHnqCgiwjtPGdONelh7jKffPVyyweL9UO27lanzRpiYikLc
iUiUm4TiCXXTrZR+QmeOD3zVXscjaSxcnAQQyIAtPLeYWZA+1GZ05Notgef0fulEIEamz9VV1jMr
EsiZtQQraDu4OFhBx2dZe4MDh3U4/SDN+Vw0AT9E77QdV+Yvzi7VYbZojCd0+X815MgWLi6RNzfW
zeYPd21HSaKBjvzRcUf5YIOisFfuGpN6ZKmPS/piqC+0BtFvtTefjbROcFFUkjddGocqt39gloYb
Y8L2vL9OrS4EKt68+R1i8+9QzW0By1J9YYxv23IQhSrsK5QptuFdtav4H5g+G9l/DoIkf3yhLpRM
WpDGIa6prpdc3Ttu2JwAUPf30RsFfV0MjN7rXlAOtdl9YGML4nwdbP9wXFZ5brR/BvoI6JTHj6uD
UKE6cxDs3Lgfr3yz3bw/XQo8Bm422kl81eYQDBdcAqcWl50s4v/C1EpRqdUqAI43cJfZdLTBMOSO
5oowm4fL6sJeG8bLGuruvfLh6wqTJiconKBvZckhARYikWdhqIQYTF5fbJNczK18Cfxa9WwpgYXj
VGVjZJh/KgQbjwktrqBK2jAPUYYgWNd/eBU1yewjxssUjsPbce7CVXaNjrQQbqvW/7XQ0SCTD+2L
bOosmMymc6GNaSkHaEK6Ehu4+1/DAhzCpSMXMyBVwoZTfj/g6GEJfGoYTlBFAthp/zUsF+t6gJOi
FASsui4cUw4bMbM7F9/z7cYsDBeunUs6a+1tXb4GZ50TB6qTjQnfPOIjgctVCqq1aPcKW7FJ7lZX
kf7DOf+OeG8ygUM4gYNfB03RYxkqEZiGM+cfwDlwU8BVgJzKzMQ5P5I6EtxMg9aG6XnkncDg2WOf
jaQEhjnCfAfEENOOceBfKX7/M1baUVMFOsXoHctoby/zcLJtjsJ7ITL+O+rrT7fqyXI8zuMNkDpg
SWwck+NvarL6V9zyQwI05nEBK8CB5+8rh3UGa3twDqDg4BWT7GzfGXErvdgF+WyaA6FUTPogL2M0
WvBae+j4LHDJe/CcXPxXdh1Q4gL6sd81HC3sBl+tFZ3vKv3L7k0Azgt7n6kohx2KwMdjdaiPWvsy
y4Y/R/lDoBsrV2dR1Gx4H6Hva6j1egkfIixAQ7Rzdb7Jj7vqh/VIht+Ip5byJGhBL0l/QXUIrLo5
C1q6PI9Z3kUFRrkNpJQcRLKQK35JBbApuAtH6uFWVJyHgLj65SAzlfVuQCzaAl3bSlPWoUAbTWTE
WOiiGq7m1tMGmg35fQbNgDgZ/iU/ApvyvW0ANvZfA4RI6ThzVA7eG0OvE8NrPrS6+gXuM5ASbME/
cTLwqK7ZsMl0qCNLCF5KAyNo9V+6ZAHPMW7qoVOaoDmw5N0qvyxA5bGG3YByllb/1k/zQvTD2EXD
UhF6qPqgVe6610lcIhiaAti8Jm8Zn7yF9LEIQyerO/7eVozd0uSlDVRFRCsZRvE37yTMihAUozFn
X/f9wJX55UvK/vkbKBEKTSqv6YaCiDpol8zu7R4aDSiwPm/v0gl2JzIz0ARv7Ekdmh7VRtr/jkEu
dyaoUGv7iDGI+HNAnnkjVXp0Ila/SEnu4eGj+l7U1DMzbR4fQZkq7sSCGNpdN90al2X2F0wIkm5W
x0rRt3Fn1kTRvI/3xauP35ZPBUMFHPwpYmM/G7jO3ndtHNqTX6GfObYxT+lsvy7FwNT/4Ixrrygf
toEYzO5tWfuUUuuOtdbQwEQh700TptvOZ2b8W7SZCEQYJ9gv2SWEe9bJ1E7WfRY6X9zkgA2HmqMw
BnzPatJasDvEKLoR3IkJDTt4xTB0VRMoSPuMu9QHgTtVBO+Q1V+p+NEISsDnSsHOjH/ajQAIJNgA
4i978DRMFFdjZIghHfiyjL1YBBn+Th/x3aAp/bnSiY9JOWXHaMjOVJlmX7V3hWd4kka2SQ2veg78
375z/6TIaEdLIhRFW9pVXUUsWa3xLpPVzbozANMxZZ8+nHwtD4IM+Y0O0gBDQ+BRrDyC5RsXEjvS
ZgLpUKh6XqL65oOfTvyl9/ivvAxX2JYqB2Aj+lBu6YSGE9scOs6zXmYyjD8Rzm9SPMA743qgXGWb
Yx/DnWguGh/x7VfhKvLLS5ZB3gDihAsfVaUxG0crpQU9aeUXOQYgaUO0ux18k/TlRHZ5YLlzCBYB
uf9k/FtiMG8rsUXWRFuf5sOhzwQ1KdP9tv/ewRvGgJYbc/er9pEEux4jNb3zMOAErjC2L/pAR2ka
bST6rDAFqh9gxOSDHd3LsDC0T2QK+XMRpmNm/ahvo9x+R4gXuEiEkp0MaadEjHMPyd6zpPOHf+xj
nnfHIT/vrKAEX4coWrZlqxyN/e8CNKxtxnrzDt04PzUiGoC7+32idqld2YZwS1PSEKjohCY9sV/H
YSi9C8It11STZbIePcn07kpl4a3PZC6CgpivFMHBk7PO4dMMgsnTCE0YMHEi6isK7E1EHjFAlyeN
8bxnnQUvcSoj1mwesJQ7I0Lq3v2QhRuc7NYadJa/bwhNEUakGK21vdIjcvev/IiSJef8fL0Ba7dB
mv3netMbXTVwRzTcPZohOGkKgZ7ckJKG89+Qmszui4PjGBrLA82qD4J8jw+axx1sLY+dRwq2o5r1
hJikWa8YKHmeMNo5Y/Yg6GOvrlSuQvJd7dzDjAbycJFy2Uw4KhcuYbKJiQsJ6VBswwYSGTdOa+bo
0PxgSpjB879IXKCc/VSxwfxmurjS3GossTC0oMaOIMaRmfOQ+Da5xpZrt/sDMQDE9Kzmioji8z8B
olFKCIkLQFTXQ2YpZ9XEf1CQcRz8lSqsUy+37uT5WkR0wMpRXNBWw3U7uQ5MeJEwsiPdFhOw0xv0
QqbvGUydbOM5aNAAxhrXd//e6Jruqv+udtAQytLnupvsYDT0G2/09MlAjmArl1slGUcVx1P0Jro1
K4yRM8BA/emSv+AodFGVk5jWspfoLhjRzLSP3zjBGBvvSNMPVJXImyark6gZfraRVj6V5twwIy+o
L47rvAVmTDJjFOgs3Oqi9HRKkuns7ofct7ZMYKI/a4+bwy5z076tPi00Y45SC+mj0bOx2hyt20f7
bSxPv8Ei6/WfN/qKL4C6mgoPIWqAgoEuSTRwznkjH/rDrxatdSdSZWGKFYcvlVsyjWvFZS92ffDl
hwkOYrQgpj2cOD75cBMdLO5XjA2NpHe7RW4qNYy8+Ts6plt+018CaizrwdEzQS81cgZ9p7Gppzie
HwM27+tWfoOqwWN5GTfAH0tz+EDZriX+wDYLqRT+QEKxX2gJ6Lg3ZJ36+vgOKjaFwEMVN9/sDd8y
3WzY9Na4Vk3CilGxRFcceXmYr3weTh59DaPQPHDWYtNhCihmCGANXzO10bEt78jAibvMMcZWoRwV
Dmk1eTJvZXGS32e88S6RZIuxX+iIZbeElOdEE2pEqGt7CSFmEDMGSh2RChPVEoHXgu4QuDzNpVjS
9nC41ITF3nkWx+J0cRfXfLjJzH8PaBdefMurx5fV6V4T/9Q4C3EM8NYzadtEYMcNSPnfnD0V4vaq
yb6TA/EVhMa4K60201Z84/DZGRCJAhYf8/hrHcRrtCzVJGDdLB6lyYS7r98DVT8Y23u1NKrL81DA
3wXhMLerS6qYv7bCFWs6supLu7e4YVxQSfNS8VwKlRuZAh1vvHzeeqMryMTcfNgDvgAP8Xrr1xyz
nMOy0JpboFDyMK/+5y3GKwTILGS3bWWjDBi+NqUMr7xPfoMIlLRfqX2HvDkP0q0VSo0+ziDaogRl
Ic+F3/GOFJQKYDRMdInHHfq/lCHQvnSE0O53Es6Sxn3/10tP+OC1pnqs7zYw5x61hhtv+BY7fVD1
r+/XxO93OkIpUNHBoDeV4/7NTnjs0WG6ubNPcL7PVwPgyu9dIjbPFwjXWEiVQZIyb8meGLZA9KuE
b+uj7W/+J5lFDZ7ArW7iboNvSwcNUvBG3YYn3YFD5P7aet//hMlswBizTt0tzCi97s9pCb7qUmiD
KEWsP6PsrYGMiDRcCrzr5E7T8rXIX5X2NVWnWesCD0NCOg/y/B8bHfkhfqE2qFtkhj3nClxuGg4M
NSawejYVhb2BS45Owtw/6GHTZbO9qkkWUoh8GyoFCYV7GR+UAtFuCuIxCu28o2T57Zs18me25Y0z
XsHF4oH2HOzIPKlizc4S0zWhRY5enbchQsLK5eYjVidlm3J2VKRxKr3Uz8KgM5m9a8isjE/5xiJi
4V71ef8z36Kg5Ojf42oBYFl0WjfqQylNmzY+ISii52MOqYuqoOr5E1MDDQx/Fw1AryjtrUBZ7CIg
7P3tK0u+RHo+eQYujd014O/D3AnQP3KvUfbn1Hp7Go4CPhqRSD7GlpYhbiPTYGyfH/9yVWDbDNew
9kwKX1E/O02HLcjc9D/AtoWEffLBvNYBv5BehLchycTiAVW89om+3ICVEYtCYRAVake4zqjEQlfr
c0ABqQjJpCKvJJYtxGgpuS0EHABTn2WDrcEB7JkbsG1LRCXGImvYIgE+iT+2pmqna0eEKDWEaVA3
8B6F+fMFCzs+eL2+tisDIQ5I3tVSgzSKvRB7w0iLRubMKaiZZ8RL91ZMwgvM++zgsgXkLousXeGY
dHQTFIlthvEiDfTRVUy9E7YFCmJKFhqr/x5qEFm9RlZpYMS+7YmmU7xFWMNUa2likheKEvKfHgcH
qst4DdhvZ8TfK6Bbxavc2pK5rWLsllGnufRQXCdb07D7hC3EXrkVxduSjnuoZRK5FfwRcQgkwb7E
gkZ727lvsGouEYP3R+N8SAag43DRFSF7fj1nSzTtrvAZ0+7Kmu9MNXIG1R3nxw+Y+OhxAefeduLT
JyKIWumkx/reZ7b4BHNbt38BCyYNXIn3SbZeO+M6Q26F3cV+qyZC1jxu0NTUyyXXwTgvUDXIsFNV
LclKJ7SK/9GB+GFMfWZ5gpvxJw+7lWIjL8OwBcL6wWLgPUIyAMgy/n1Kb+ZkXGmTNOFnkEW4PxSx
Zvt3yK3MoW2uNH2CcRKujbuSp3dsa/gp4xLO8fGrNu/jcirnsa8on8ox81XbvjKT1TJKcLsOt5ka
7S/TlIuTpe14qsxVF+jg49CRLMPJZoFtkOyeHVzoHPxj5RldYuL84DtyTy81b1IrBHZnia0gcF95
dCJrvaCVcUK/595dalMy1xMpacaN5SrGsNx/VU1Desc8fi6WBcuae9nnfCAFUB0+XFXmwvicSOcJ
HMYRKb/aOL/wofyb6mMDo6R1oxMaD7JoZh8dI+BY+yO2v1VZPjOf/tZOJZn24tzeETsc/5WjsvA/
6DtMqx6uGwmWViD8BWvdjbota8WwPNF5Dx4RZELKOfFQfxS/YDRq4+on8Tv5SeEYYWj8l+dc9aKb
o1roLDeHq7fXkERvIXj51QXnBq3jDD9yD1SAWaaTJdDj2dEzN55+v402dUiuInvdmrxpFIUvqQH3
9uiQQOaYdbb5TjXNlHm/2+eehRBFj4xtYJqhLeJu7NRuxIVOZdOBHvo/LlzjecvGUW3bhxp/ofRP
T0D+QfDI/024N1PYUv4bl82kIeDZFm11IF9UnadzV778IQy2WKRUU8WQYJsk8sR5+jYlc1vwUmqO
xcY/E5w9on5amoo5X9eaGqwwa6rWKFknlch5pUlGVGHndm+nVM8GnhkH8z3DNcnnyfW3L6HEJ0NG
M0WciPorHZC75qg4akzye0kmjdGPfZ4MSS5YVyBe2P/QrdtDP+Y6nI1ffNZkN5WozqvzFNTTjpMF
n21Iy0uMhwbagKT8LeVwNUfvPmsidG1Rdw0yTahIJ3j+Q5cnwxXqFeMtLDMuQG03Bbdc6BhfaWB/
bmsEykQiV+4xdn+lOPX68hEVgRAsqSWKQ8DfzVH4DJJFVmU154fJibuombgNnFWXQtS1eBeLYelu
QgOgVSwBFhkAtdPu0pdkdroOZixmkSpLKVZCURtE40kFztDycObkv2C6yaM0lhJR516xrxs2Fd+n
XdClyNM88LkHwST9sR3BdhKFxHhN0Ops4JvRmidjuhSktreBMX+PxMeYLwDcYngU4lkfiRse43nf
S1bZ+wuUf+OgOasgo9RnDlzM/z6c1x6JUZ8MIaWWo+6WNzMY4V1I1epv4KTLnjSUUFOowRKIhHgA
fC5+Fmbeec61O0CtSWQNR/HM3NZmxdMQGdWr8Pq/29Wq4Nsprq4s0q/aCn3CvMAUvKu3tcWfr30R
B9wptVzk7QuriIDz26KKMgEHGU8mXYWlXGiU+QC07KnqGwZjyRW4r+MD+YrAq5LSPwZYNH7Uk4aE
EuWa5ab6FUL2MnKL8WB5edq1vmxRg5q7RIMpZ81ZFPEfyX9DFfuQjOBP3zLSTkmO4lfsUr5Q4ODU
YochzBwunpHPy4X/fk4Lu/Wa4vLAg/8g0AdTvk5keLFAAyXOYwzRHJNGJ74ZQXneKhtcudIwuZYV
xh4HpiLvweET4FvfjNHrISY5Xk+9+k8K77Vrj98M4CzZqJ0PksfZ4z45TYayuPymtkSDM/bkG4iX
U0ZeQv5/tW/D8wsQ51EP1+B+RzOz9Gtl3SBjQp5vO29d9++ilfTHiXbn1PkmALQ8zAo/fSYAAbVe
Bosy1xL4/PlCrLtZl2o7etxCLypp86vC0jbxsEFrIkog5rjnNMbwJnjtW3hKL/3DUkBxSHv1F+EH
lyA6xxoJ386XudOVAHnlR7weAcmGeRjs5lNU6NLSOJqcCNSdTmzXcRNYLrBEW4rMZuzCNWF0cv2y
LeTkZ3nOKEsFgIaLMCBEwZXhH82x+JmSL3uD+FUL3pPYL85cyS4pPJhnooSGOS/ySHx/nj8w0ajP
E0Cu3eqjGwtFF9267M5N7Dekhdd2SiVy2wLM0Mk5EFBFTwoRtXm4ta5JqeWw5pvroa9CQdbOHvLX
kXPXoEqKR2/SW74CsbLy480w4wCLg/XwuVt+3pZcQkuJKYMANyZqJM/o0yiJ/iEi6fYh5xHTkm8g
lrgtrVKmL+wcORiT4YvdLRe8r7T6Zqx2U/a+Z3GM5ylEBACNBx/qg6L9jgMQ9UzJAhOgAI/AK9mo
yuOxok7+yHYwRqa/JjJ57CQD9NtRTydul+48DqDNIdnSwPtw9E4SAqbyybcBavRsBlw+h4IirOMk
eVyyTPHK4BoxjqZcTbUhJtRoQseYYZ/nrsK8MdLXB3/yiFc8A/FZWrsceZbit5EC7ocYC9IBzV3i
1YpG4yfTZwAimJ5rhFag7Yi8uhgU/6GcFXo93icGDI05CSshZyXYLxAUOS86XaxPNsWgFzBbUGfG
rE+T6xKLf7YaNqNRsKGv1mNV8xyf4IslHwoqjP7Cb8HCGCsSTVRY+1ADXTipQPwcCEPdUmP6n1mM
R5QsWVFjsiwJ5Z1/f4mJ9CEGEOsJbItlSrSxxAnlcrEcVV/4EO+x/QgT1GxSTW89w/sixu/0n8pD
OyHf5UkyIrhNlfBMxyib0gy9UO6dEUHKiS8k7iG31vNoFQ9ZwpPbWYqW8zC9tHN8wFtWcS7Cn7v4
9Q2zQZBm6pQQXn0utqCitg8hoHg145gXkcennAaMVIMxV3rVLjlOHgAgvsYqOFwUEw2FlrVdoZm5
/BBJH9zFBygXCJx8iB0lKq3H79i/BspJ1hJATM9Kmq6Vi0zKYe0/QvyExiE8qMHzOAZwHPe09iEW
ok9TBMn2SGe1PUwCTEeTjZKxv5COB5J2J9sHq3yJ+BNzo1GExiGrjD1g4JO/6JexfZ0jOa00gDY1
g6cgNk5BLUzPAnLbCQVo3RSXc+ipKDOalcxFlS3kfk7OGvTtKwmpa38P+7ToJKgUcLI6b1u6CH2V
Xwpbi1uBpTEiCwdpV2pRyxrDRtu2EJoyQ6whnl+cOZ3EpoMwUlid6ZBTVW0/fPB8OG43u2ySFIKd
ZDtNjRDJIQj2AQN6kbOzfyFc2qzupMBZV61EeZQlaks5Gc842kWVaTNxzoGvGrlCHifWsFKPpXKA
jRAi6EzG+wJH26tONfWqaS1/9XEB/nSUVVbJRB0YkBMdlHqV0T5WYwBOXugBBidDtKd0sbTmVZll
qlVJ/Z4sb9FCyfZ/YUYsC+O4AIlY/2lzxbT6Ya2IekJRX0NtNauo0jO6uNbgyKLuOhnRJ4QAyfoF
xxJ9OKnSSuxCq95kvhYgQUuDuYQd/MIJPp9hXJOAW692H5+dVIs9XTzu3PJ131uQu3UIHMGxMq8C
dSb73B9IWWZ2wnAd8WRLd0zmcTwIdwNq1M11B7cj3E9anWBVzKI0hph0Ivp9J9aI0LFnDkk/W9rh
CAWW+Ti2jIXFHwbqVbjKPJmu+WB6sdGp211bIHb1/XZdKlg4Y3/97VusDW7jA3xx00GWyd0oWmyG
16zJLLWFkMiNdWTclgA7PCrDsqscdvdukJvgwSw7EvDJEbXRhYengkfvty8raIs6NKpCEIRzhuS7
gBV/ezUjjciVNEiFjGzw3d9rwKDvKF0sez0hLF8hcQAKBUHGtaEM6ibphI6L38qTKVUnAxesOs8H
en7xnANvgn4gtOpaUH5FbDrnglmmgPIr0ZCgTLm5HuRxJi0D1yC7zppJjj/QxIy3Iu7ciWL5V1Qt
uOMrsPLD4P2uQvLuJ8ay8i4XQzIjkUSiCs9aGqu2bx864MJjdPzIa8KGBbnGih0PQfg6bThiYV2X
xIKGU+O6nVTNf6Yj3r5DfH4B0J1Os2uWSR/DLYDbXxcdMPCiJAV/6zdkawJ9FiSnxn1Kavfq7EY8
Ze43ypYDkExhQ79fpSJHfwhjnolgnkEm20f8b3OU99Nsd17g0TsBCwyc7j3oUxqSOwZ4Ay1tbEI6
Lr12raWW2aoGD2Hcy30FuNFzsUvntFq/jgdw6EvqR6M6/tODGz3OhaTDyzZtGGn/e/wAm81RqcW9
GIXjplMy/G7442oTKYm7QKBwEKXwxTYIgod+opLdWQvWQYW8/IBdRRRcc/0nRHrQjsAj/orVUKJq
ZuNpjGL0+evb+r4hSh7U1dfo4gBFGXBIuhzKqX5Zep4bUBOsB/+Nqzz96t6WgztfbIuixmeEOc0D
k3H108fGV1hdfitIMhnByEKSwMXNPThUBJoowpJxTLo/qrx3qp795V+hil5HIxDYWoLmI0GlyQV4
G8cmTLWztq1cm3AaJwsXdlviXSBN2uzsIAWLBZPA2FBP115fxGiwHn1lfjsUO2CFZLoaZeVJXtx7
Uw/LE1Ruhh7sOjz3oNXZxZ3HvphvTgVezVMgjlcF7kCIw64nxTze7LIiAp4xuoV0keZHuEF3PY7p
sOMtPQ0+DAvXGiv1aXIiGBvKs4SJtGnP0FqZ8Ur7xHO7EK8seP5Sr99BDXCXuty7fcZqmUZKyyjZ
ko/KvHNbFhyi4JItkLHuojqxqWUSbx71LPBZwA+Avf/3vsMumtOUxeJLRX/kOsd/HzhjAZQkK/Lc
VEg8a03Ap+jVbnQmIjeLNAMQjoWWi+KKCEaAHcskHwNLlVyw75re73KYIGG2dMrA4rHuyRdG9iut
nzh0QscI7MvDK+w4mpDJBJ2Ev5s12MUl2BbOXtltk7NHC3DyBv1rVvW37VCcCcNud324B+n+apay
zrwzNGSXzYN7RiUxgYvdZ4wLqDCNrnrhTDR7lgJMCqkt0VoqX5FQ4Zt/KFLmHzBht840RUFIFFdt
XJO8/ydG76/v+itVUuhQzNsAyUCc79PC3HycO4az6ZxuRPDaDA54pL84bNfdRPDlC3CNzkwc9vR0
+Nw3Fa0Hi81tFMfDjnF/tWX4MKCJEwgI7iPgwNR0vufvGsaTrPwvnakWdYbnK/8t0Pn8TV4VJeL8
pYkLNDu0yAbQU7Y0OwElRHv2AGmsKJzgG/h/ok6RP+sH/DaFx8S/hMexyng55E/irU4hAMzxAvru
BvtHug71RxwdWrWQUFanaJO8brVVYFiwBQeuAaUhu1Sm3DrYxP8ppdLedXVPF2sMD4EoJNKqpcnr
WTZ1EHWGFTR7MHLBYUC9tZ8lxphwRCWVV0cX2X8hO0byt8lweXrk7WLM/2swmkMWDyMHKZVTW7VA
x+yzXHPr5jzTweazRE03C15Ku4UYG3UB9MEa21YymJpRqw1pnCh8tHg/zQSPRGPsqhpMV/ixdKD0
Psmu+O8/vr5k2dgPKxzYMBqm2Xe9pUgM43Hf10zM05NbeL92w6uRiSksC1r+y+M69NkV9e3c4k5m
IVJEXxfD7povj7sDjGIkGDJHFOof4lampwr+1T21qJiwi35CBnZwAJHEEz2cKLGPdyldGrNUpW5E
rc/GhFdAY+V91MgjQJKAc6gVb17u1kh50ElMZpI3LpQ+q8cxDR22KBQwBeh1V06ucrhRS3GDQbRw
dO7djDjK3k3I7+Q4OfNmDi/AzpN1K3VEYL0tYBv8a4W93cASCYbhGF7nQCi6F7/qnO5W13jmV9cz
mT+S8Ztc1bUNh2oHkTf8E15UT5vlq5zW+uHdS0PqH6g292T8mJnylbjl7CVGsyojM6iRyYTX0VqY
ezWYH2kvrghu8NVg+/g43mq0sfHPtjlE7OCg8z/iHxu3RcudYHQwwWmiyvjDHfDKAyv/v9n2T65n
0j78DnJ+A0PEBDkgydTdHUKHye1u9UiTD11Nu5+d/BdmK1B8S3fyn35/SgA+V22SpGaMXq1AUTZ2
wZv5j9L+/NmQfPSpxDeHTnsGSfLmBP24ASAlauxNfkWGNr7Y3G8hPZ9PJMiNT2sPGj2UeEhvE0kL
DINV3TjyBb5JKP4vizgQEdvqHxUYQH6jc88yXK2BquIt6fHX+jckzy9nd7N7ICioNNyP0rDdWsx8
zqS7/cqbHUuDf0dfZj1AldyaP7ZEZv8s0WH45OC51a9dr1XNwGEyav/dpgTHAj5iMd+Ay46QtzlL
GiRzeHE1EraUGPY4WbM6xZ1KL5DTNo/rNfge2B2Oxp9HeC1S7g/GF3Zxm0XamJjj5yrb971MGjcG
wtHGXTTD9GrSWRvFFGv4mn5oUVZ1zCyHSLeY8o8lmpafRExyrZOGP1YkYVV++YblQU/oaw63F1oQ
C0whf95LC7YcP85BHs0gwChgVMKph/U0bEOZpaquNY4MVmIspATTqWrxMRLhuv2S6Z2tq48PGea7
QTzfobQvJnAG37fEx4h2/yQBqQtx5mer7N4CdciD0fVUi049MYjhtEWwmGj8H+Rie0R+VE9ztHbt
r9sz6YAntTcX5mATVg95uYbcszOSmAuMTorx4kOL38N03rSEtkcI7XqmwE4V6sJo42qlKVBcGebi
OU7um/7FZnm8sv9eHXSKGCDwvp8VSpxMwLTojZGOp+H1/5kbzujncPwp7+FZlYzFJmjGMjrhwjRM
+B8yws7dElv9PqioepY7RwDusM7uHbbVC9H4mmPU9pb/QbbrrZeSPPsF64qvvxuMulAXEgdgCgK8
V5pxJdwKI/jV/qB4Kt2SR7tB2q5M5iA4mUWTEJCKVY+06zlOXjcu4GCuOTV+kTmeYEde8DezCQas
i4J1uK9H6seOiz71aHU1d19VjwIGWUvS0l1Z0zi5IpT85RUWkRM5PbahLKa0DmgIBcJxWf7HelIs
vnc8F706mucoV9cpb3JJRYRf7QD4A0hBgriPwR2Cjd4Q3Y9P8FcDWpS+bvi3LhVe7VmyoghwjpoG
yJkN2LJ9WHwb+fHWWnVFZiyrFw/55Iutk56wxzyc5/XelV/NS1NY3sdmpYyeh0cPihF1zFChno+7
oVmVszaIAS0xrdt6q43m1co66OestPLO5M418zEqShcA62sFnzMVF/NcX3B8gUxFWAvrIzlwdNW8
wlfwXDssV95YZHA18bh8G4iwAKfNOFwdIwkzPNcQkKMKm/hZLNsOyZfmGEioM+QxwnYagdAOmHuG
iDjfjedMeMMn8KCfPI2r+4NNtrOpFZhnsRQFYbG7WxE4VeYG7TYuK3Xdh2YD/AhG2LusnqZhJ8JR
nRE+b8d/hdawiFTkdS/gd2PI30JcTY5JHQsVw+28QQcF3WxQ9Wq+50ypdgAXI5YdjH9MYO6oSlge
zBYyHvrsTH4A7PPv+BRYFqEPYRUcPOP97/gvQmGKFP28pymTiHkTAZTPj0uzSG/RfMIX28grAXw8
oNgiN0PbHBfUL4Pnk9acc1fRI2mpX5bdHPG5VhAx/6P3Lt+YxFVvj8fwU34SKjk8JtZMp3N/t4na
4cLGaZT7SKNN2cs3AN82L7x2cDBQTIxkztD9C1lvPi5erVGngZDxXChiG9mwvDg7UekpEo7W0Phk
qZ6N2eFH7JAhkPpvlV1id/K6EUKhIZoTV8W1N05x1Epd7EPKXOJiWzKqCExfpwRbsaAbDMhZPM2D
qxEBqalDc5MAqxEs5kayQihA0HncOxosjPTpIcOaP6TUiy1zkfag68p9l7Rbl8+MMPXdj1J1e1PS
YCdXircv3tdkx8N7SIAJfPkAZXyzsCk2Ueo0CzMFA04rSNzU/VorbUvZ86urIgK0B+bYDLFANqfn
KdU74hTyhr88P5tLmubyqL4aJzeKSjARZN1YjdQ9GdB1qRw1Zbu76UrMsi7sJUiucR39bnGoKC1v
Vy1ZSfJjf1kb+o/XXyuxNF/KPYAT3bfMfzIpbd0g7BkoKQXL0BvbumnvT7TJpjg/Z2Xy3SwO9QBX
h0xSTeERCrqtEZ0g8xlEL5U3ADkDHFlT9YWAinNmo+Vy1VOgO1+tiw6lKybCs+RLPTV1Q71woryl
V724FdJn00Kkd1IU9g8R66ntjyE9YsFrWWJ60YMGGf9+JSfjb8PP8FDJSJKGt6vqxPJw1OTT48X/
B2TqC0L71YWygIi9kmm2CyVbVMR0xgkRnTxEJjT0pWkf+ROnMqqQ8Q6fGQJ3G6e9D7FjSPpB8IhK
M5kWgLt36IjvNXexJTHMKk3QNpjFmo2deXP0Ng6BUK4j8DLpMVeHclzvnNQNBE5q2EWum3BJmWn6
P3vr+eL6y70A7np0GdE8I76xRZAMtfrntKWVlN3DTU+hVf/DQj1JlmkI4/MbtMcmJz0LdDtEXZ1d
8Am0bJX6BrF68po/cysg+nNqgcQ7j3uMfEWTHKbjTKotKdp92l9rniAJQmSQcpsRyYe5vDFB8t/3
ZI9QLad7+QCjpuYKpFET+R+MdyQSg8YG/kWnCps0wRCImDf0gWHRYlCesQXchPFdOQD8140fNGeW
geJMtu4WH7RAnMZYgfV68MITyOz1QB2t0Cr3SKCSVddnsCdSrIVwNCtXtOe8PeqULvjgAcC49lRy
vKDJkuwweIUuDWAlT6vlGs6NfcCTidTyaH0/0KSpLWXEeQRibnmocQ7VdGst22FSwB6AcAlsssqT
ML9GY4LWIAoZMmtg+uVaVELShAiDTuHPsoqXrE5Ymrx+RimS1VS9VwDU0feqCZhtd1Xy/qkLx7Aj
P7EgjjD9Xp0+0qEnWdwenYmC1tSJSuK/AVfgDDEoIGLv8nLpUueOdMgSCEsiWr4ah/cm6UmLqHeO
7fb05WOWqmCDdWPoVL+bCHPGavQtMZebD3N0sd1x1Hg5h7JflUNTEfOd6NeOLN1TX5O28aL0DSHd
O17kjtKrzDxXYQUdTmtwNbtsDDgRkPX4IUDadLvbibvMGzVAVd2FZ15q/jD1L25InvJlLvIf7EQU
mhwG0jngtX1ejpdx73gJkHTssDQoJ9P6LScti1rTAqL2k64NN1D8ipEbWW7xaZBmZzRXfPY7TnlC
HDaUmc1XGgq1b44Rlg/tHkpet0f6cy1OELDdGoYugSYM5iQhHpmC8SBo0hVZW/qjGnPoMAoDDA+B
LDj7R38obAElXXbS0oAIaxE6/HTcfWQs7LRzEIucPTcyFbmVLAU5R0yYUACsini34J8ESrFwgaXc
mxO5GiIH8A2Bcnynpo1hb1GqQXMdNSn8xQGbvOXCPlDgiDJXe0We1xlfnf03KmyrZU9Ou3ItmUXV
vYDSq+eplgTPzIUEj+vKA8CdjvIGnTA4J4NGQNmJI8EFAV823lQVdwFdmKU9CwL0ItEVphcs/MTO
qbzNqiNEpwjI+4TFwYVZuA4oRH4hEiZHt+lcWOrLuwMnnNFkz7FwVGfVvyQL3YXCYdiWZGxQPFs+
vGMRxvFjpOzWoESIJhHbXiqMnIQIGLV7T5vgpPRhmcoJdS9lRtEgf3b3yR1Pdm9VQuagVcuwtep6
8win/i8qwyEwjb2fUDVqqxyYHki15wCv95U4B1aMjHbwWvVOp+TPhWeqhnQNMzTm5FtJKkHmoJdM
WhizLVTCraaOaCoWDrxGyF3yEPMUfx/T/McTE2Dpv77yZubL+j//ILI8QFkJk7H6jO9j5Uul5X8p
3HkXUXILu65f/gelKKbYDnuQox13YVgymJtOPfp991lU7ti/1VItzYLWeurGQUy9wHDu4IpJg+x4
GCKIy4mb31lwSK4MQ/qClmGJh5kCy22dxNgWDboNZrNyOAkKCQfRxxOHxLc86kvVSOcxWfWVsJN/
wV6gixLpnQqTKWbGL9S6fByDyxkpakHYwyw6vnyiYKea6FlR8by9oVRjr9G5X3R46HkoxrUbb3z/
bVdCHKa9/P4ru3qCO4VlZGIEiIvNaJupGtnuWZ+KSKBcAAd1S459yFTCYFHQlEIlis+cFNQ4iMFW
UYunFVlh4XmjdsrUWRgMDsWkrcxr3hAxPQ0o5Lz2Mvy2hvNgwnz484XJTbBRPmBa6BdtP8LDa44q
sT6MbCCiUqHopp0E+JdQuhwiktjdNqEJUuKkdC7bwtwsfUnvlT/zrpPVLPQtdlc7FZ69oTjYtcLE
ujeKuaKnZN5BSf81zonasLwSGg1wsYKQanU8uG6RL7HV5wz31hJ4uApaZQbakAhgnKnWSLSE6zyZ
czhqealo2auJn3a4QPRNo+s9FH+Jw6uy3URGgtUxAf5ECxWFKWzRR4z7IZw5rX4N3sf0e9qSKqgZ
VfFy2sLwODSoG5gXfRH5tON3TVhKNFvCu2/RqW0hZbCZSCsv132JBikxXGL33nRhPvHA6h5KfXf4
vgKkRgL1wHNkS+O6GrxI/Yy+10sQxwfC8i7Y9G/4GWvZ84DNNhW48FSUsqw9zvCz1eBBgTEfXfPq
mtuzImBUbb9yWlKpHhtVJopPDkKhVAr9GZk5FQRr43g4tg2QsRVHnhHgJtczpaQgzTc+Gs88IkfZ
YXcMq19dkrhOpYmlmlqZzbSif1Mzh1bMyY/O5CngtG1VDyuqbITjgKAP1LdsqnUphIyn6mM4GlvX
gl5LozXoIw940XLwkrT8rgq6G0B23Lo5Juz8V0wsVJfuZoMIdsiuvN6BeVX81znTplzQJ0L1zIjG
uml8QLSSoX7xhdw78OsK3yDNqe52s3ycm+yOqTOnmxx0UkFgYk/d7S+pLKGvg7UlumHRZtHHLdH/
m27YpUecR3IUbuzvc7C1kuohg4BHUkzSsC/+K8tb7zR6wqw4tzclgLjVoE8TJ0XCHvizz3cnkpL7
VOohlCKTW8BdKdjSjV6pk3q4N4WwEOD/RvGV78E9BnERSQZjSZD0aXZuOyvqJZzkrF+AKYqjtFa1
iHzoAqA2qo7DacIHfpPM7QSf1RldF0SPp528DmOxwsGJ8idzEhwsFRRs+l1O7q7rpt0jggfpnwDo
A8as1jlWnO5S2oiNM3NRQqZ+53VaHhMj3eoi0tQTiTttK8ZKq4klbQSdDr0yvdKJbpOk1zUcc48I
h1wyp5ZuHAIoDG8ayzpO/H8U+YlNoz4I7qL0FgQNDroBPAeZv8dJwyNbD9RAf+WON6OAV7hO06Ab
wVktCLl/6G5Y26MEFs2WiZeZsguL2rSEB+ZpDzt1xJIkq3qwOnx31z41qkg8Mf5N/X6Jn+uATCo8
Y6VHa2beYTwWfRObsWYrF5M5eu/hr/t1NlN/qFQDl30NvKdioS5WX/Fgd2tt4KRj/AEvMmXMjXNI
MBMMfElIssPHR0DIhN42wAotYBRx/tUlDilC/MHvCI4PTCFlTwV9H4JSg4j+2v9MfEva37lV5r6Y
EEpLUtDkBuqs2VVQrussXBibDblZW0qOdD9Gpxh9De6AombjMrESAHjnpB6GdFxKehjI83kwKm/n
ZWuxijl5sdVknhclmjfC/Xjh91YE0113l/wWMqgACLjEma7EcfGfoELrcdBZ6Y2eoGi3oC7KdG8g
4X+1ysuIOfFdnfTrQWrKawOCEVDxz8n37axh7vGsiVjdMvmmbTXtieXLKJ7OOn3Pl+WNGrghX7qK
K2P2ycFiquxFafq4KZ34++526436ml+4/4+nDTXx1j8PetKx39cq3K6ypDE1f6fh6HxeLNWaoDne
V7g9MlK/YdA/C44axyiXE2ryM26XUkoY8iaaP6Kf3WG908MenhfnrRCBkS/jr17fCChzkTUUiqEx
m7l/Hxkv0TeM54mUWDv7kIw1mtO8SY8Jm54V9FUtWkhy9NfctoLmMOqBX89o142mQgh5YYMTknz6
LFWgn5GfdQZmpqBbT4JYWuAqCL8pK23xyO6/ReqEprbO8nnsLNcEitros9sz4C2te0JJGUfk6S1i
wf8afIr2pOJ5kr7636ief5GaElVCY5wwFGBAo0v6hQLQolDbkC0gkTEPMUnXV4HiiCCgUUCTYnh+
BzvpB8qKne7vP5YIuhpvVFX4i32eC30u0FoR4rEnQg6dqFYDpznkS3E8E21atVIs+5Jm8letMdMC
gQyazy11OzR4rtY7YDMYuqrDT3g+0NnQoPPH/nmDWNIx0jYaTx+yxRbfb+7Fn04ngNm8E7aIyDu8
n4T7G7cv/7mhA5v1LP4TMuw7xc8KkYnnjtuA2oda4jlNX6lQY6iNoCM02fZZP+gYxqk8I5y6vUFL
2uzu0bFPWLKdmNQgDwuiLtf5XpnajEOgunHMkIr52FXeRdw5HipKUXYfXl+STROUBjFMhhr1Vi7U
XIOUkYPWcv0Rfcb9VImy7NlsjQrY4NR39eSzX6CBag/jFTy9mGcP5Sy/CUiMC2b7J8f0DraotX4d
i5ssfe634+e23m/RwXzVmJi+OTDCand2GyS9xKgAz6iZz3itUQ7XZFXkjyYB6ZumUNVKsH/4hCQM
lmBAkXHAZdAODYct3/nEq7f6iUtC6NAx8gzarPamV48ND8YvsZz+jdEU9n64QZcNwwEqlnJqLyXo
meALoOCfIXfGasdi3z8yvfm/neTc8Yp2jvk9QbIomApWMrvy21vsBqU6hIrcLWvWLdQgE8qHgT8e
A8s6/KTKu+jUqcrDOm8EkN/oYlrl3KoCyELIth2l/NSjNV+kOQX1oIEx9IhybtNOomB+jEp/eP7f
vVhp83iPn5XwNZKv/n19WoYqveqBR2IP3Ab8WxsiW6s9LAJ+CrG9w67xPLmsNtFKrfnMKOzesDKO
ZTqB0IA2IlySwg07CI7Al2qPX5z64BhWCfJrZQeqlkAXqPqVxoa9RZP+FotfXOHlIdPH0IAM8m5k
V0oPZkhA475cp7jVa9MXLqBWJN9Ncr11vfKHmyod5SIc5OujpJS4aoZW8W8Pw6Ad0Obybc+AlBft
MFIfniDG+CyFU9A13cXsX0ND7WV+VaS9mrgq44QXNoD0H9AxseR5facLnwTB4SobVdNhDClthd6j
j0STHZ8ZJgalW/89dx3xvUSYfG3jvOfeDrrKpXnZL++KMRDTH3optllg4sO9vlohMw4mNDjy5peq
Ngx41nTwdbz4qYnBiJBcg2r0cvEgnYBXymaYW2qyepVqKVsfNhUmPEhwt18ORec6x7ONpiqWKsSi
m3jZHsmwP+hwOqiO0ZrMEiNTw3gw8VVAmGgiClrFOZaYMeYlc+6R7/gId+0KZczXWeUg1LHnI6ca
mmnLIjAVZbVUtrjVyjnQcvzd00lg62JR68+1jzRGOcDqYazvyXNc66eA8VJ430NoJZmyhiLGBUjE
vE5FWobTLPMD2vf07aCM1H4JOKI3WrLXxXaNuYm4NpwzjSyYf1mQ2ChsnC8NxfuDzLF4HupgOjnb
8QqoXt3mGkeDsBgWZF5AdJelmDSsBpAyIiU3WCUGkKoY0h/v8l1tblU9t/OHtqNe3yYTMdsqY/Ip
gnefnAMTGBuQidePygl9vwJDVRz8VhmG6SwiNafYrOqiJxqiO0moJrILey8lCBWgNKPkqIVn6e22
QjObnhMb+doqmW6LvQ/fMEcnsL8NtIQ6nXTHOm/fuLV0s8wfEmzLEfFG1/Id4ElqEXX6H8gMNK4C
icA1otCDfJ2GSdJHE4ThZtla72AbSEFiTU0MJcpN2YBzhloH+hscx2H0dNeWnAtDcjI1SKJjLxUZ
p3ejCPYi5oKXTO8BdSVhh5P1jkHDWoSry7Nux3cKBHeUUsciVWRbxeP5WUM9nq2Jt/K5uYeVtHoc
3oG60X4sdV/9V9n5etDM95eq+Hy1Z6LOSExLjBZCnyEDECfWy11PYry/mO2oCSGdd2VAQCLufzon
yuEbPbjCUodeRL4jOJ5bDfFQ6Hu0uPuqNlsuj7mDCvwTxBwqlGn7Jr1diwtdnsupsA7IWo7KHvcv
cx1e4x5tka/pb+rLz94lO59fwrRdTegWPijXSq4dU3VaRCstv9HFnUDg09rlwk6utUeFRqaV2/f/
6UnkIXpx0t1tlqynuiasW9rJUgbxFO5T5lfeE9ZlnaPNvkPn7B2GddTDmsz2lbD6OV5PVeLaM3rB
UG4xoVk3T7Mfyzi/5Qs+oStuJry+zdqO/qtaOKCbtb+M2j6YR7XXx9ckfvmY6NkoiREiVjeHDtYl
hbOImlXrPI+n2mjY7TZjM4MlWsqGrkN+5Iy2UQli2nMP8IAl+sPsKjvCaP6cqJ1AcH8D8z6EvWo3
9yEumh7YbP2zF0uin+G9Z6r7s0xqubzMsGeoGu+mWin2r6M35Sy7TG6sWYqWphoiiqQZpH7X7Hko
Hh/hiWb2RWmKeZkUqO75CD1qDDUCZlnD47ppWGztJzh8yIzd5lCYv8Mv+xmqyGjC6VTEaskU6/Vm
+Q5GGGjQJK5NKi7tXRyrql67vAn5eL/7PxE8Xi2FNnAD4y+RZdjsnuqiPULOdHa/P88Tq8fISTlM
+2L4awMkRE70m4zQDqhLsk8gX2OOGN0/gVY+SW7qND9i27T7Gbf1Eb7+pkELO84dSdNWaZITILqc
IGf2oRg9a8hD8mVPhyfUaLvJcZEzNJxA4WnXFd4QDGLgXkU19suVhgOKbs3n7LNJ903KjoHEBIy2
sHJHs0rkFnCOFgo0UjY2FiA7zbxqSYRdK0qcv2Dk1VSpw8039FLLolqIrGgVvVcfjO6CWZ9I++tK
lpmLgObzgOaUfprxjYyDwTeIe1KiaY/EPnQOGd4103O/rOE5o8XvxNHWxvief3bEZqBunzlr8m0n
v+edF4Hb/+MdU5tIK8SnRpdwgU0DW6dBM0/wGUFDtvjWeNKbJkzHtQ7+EVqzf/sMe8FI2GQ8g3/2
x6XyYi+GGNuUNofkVF0BTZ09Nrfq9pBB4G3KFIXZIJdRXzFX81L0lfk9I+FlOXGUNuOUexE5tuAX
FK9u2KgV3RTpVjTMfg0n0Q7QF1ylEZZeeOMRuXDVFdcik9b5WHpP/mHJhCT1ExnpsZeiLxVbt7m6
h/ig916vOXjvq6cUOyLBZT4wNot4zcFGVckWscRq/znk4T3C7D9GLoWIt1XBx5Vn7SvWSVeYVyEW
xypGTGpvFraoylWR6Wvl9jQMxbmMTbqdnSzkLL9SBfTFFKcpz+8/js3TcpXo7fZgtkI28LOnv3j9
gK5muPA3SoE8jyp9MYm3tni5Yzww7qtOHfcCQKgkB1tgLcg058mB3h7w2Y3Fd7J6s3/MKJGORzhI
MUPqWIY4LjDf3Sj5ys3/7GQPgMTgZuk0I0fPO0dGMPnbR6qrmQvwWiIDSp53YPoxUxjO3ZDFWy5v
0nxzBNVZZxUsulySnLKRvA32hAyl6ioY6TkAj9n1o/rPzgogFGwk1XYu+uHmuTITdORYa7qDeSC0
R/SEfw2AOj2/4jMejpbW0VGy1J9XFV3WE0ZDnDQNABQesy34RxYw1RegrT9utqdrp7NDXK6B8NwI
KVfcUax2I4ndTGiAXG+7TPu+OtmtkXOUnajBsgqldQlQ13W0u5NtF9opWCilV9p3I/i4D5eAlhJG
oetsKWDcGg3Zw2ywh1ruBDwx/MiM0eWhN+pfe8PpiFH8nr4YwPvRRh1//WIAuD2PpYw17hvL3Rsb
Vsrx3dSXGgb3Os3x97Mk6yAH04n4cJuXkFeY8wl7nVka5zjALO+3SKBY5BnW0wPXaax7vM4ctFmP
YlgQeeZ5V7PUeJWyqTWM0wshmH1ZiN/qfrwQMwh51bQ3+8Jy/kyFfwgVi44eapaTSVWoi4QP5V1m
XcUog1pU20KI1rRzzvDPryAUrxps8MShXTt533tGlGut1PkRj8AOYHlCdtxFVAw1MRfMHURYtn9/
9jMmEKeSwqSU3vMHl7nCmdSfi9kOPtZdN/KtBDOqw4h1L5b1YhseFTYSpRzr0ZHfL4HTQdfdbUG4
vDgX8l5ndhh145EwFL3EQ5DepSpRqanOzofMf2dox9RR7F/BxXEGblzt+yLC6xAQ3v2l7akYSChg
Uianbxkx/Bj9iBn5TjKbNI4PQLJdmAQ3qfKWuQUsETPK0a6RQlX8byTAThHwtFEJKOtMZw10rG9z
US656Hl9pu11SXzy2TSWB7COBAYn52yjkjNAb0grRwibfexeeCGB6Y0/Hi0C7MrQB47AXZtW5aM5
24zKv2Xvu3t3CQQ3KH/+fwsuQUpfQXZyW553TsZQK9G7TOAAxVtvk5Lnu2Vu1JkTxGmmQTEnplUo
OPc+ZoX2ISQTC12tv8ldIWFtqNWA465pf1iZnxG016Er/bSCYbYs8Pds4riHwXELcBeNFrDqCAWZ
FENvVShjBTrd7XuLI2rl8mHWDpxcAxJRRsaVCCr4gX9pO/l5gA7zGaF3KV+8CaSwZbA/7lcNLDnC
PrEzRiIWf0H0uEwEGyLtMQgI0QTRBBNYLAf6KABm0DnQ2wOF2ElDOSHRRLX2VDll8j+FaoYaKczo
AsRWQKov22EfKomhuSUO0n9ScMkyIDXUFRPfGoIIttICNpjzkCn8S76BUjwbBeC1iRsicjw71u9d
qKMyZ9/sW50JXQZHG5gSMutGJX3xlUFZ/k+YK1KdR2WdFf6XLR5PELZcaZP9F9PUQHKoEyyOe/A3
XnM5/aMd7ymsUGHrpln80ERZPRGtfJrLDB6ejqcPWb/klAmgq3fQxrh21z9FzwpDKfFLqUsagyyh
h7evkxljkRzukK0oXuJ1cWcB+lYp+Qkm4jxAlWFHXI3svBRb9Esdaw+Dp928j8ux0kcP6P+XiRzH
HALBLbyIxWp5D2AZdvY9EqR3GzH/naw/5hKkHQkN1z0aioAUFlVh0VnWpCE7lzQz/BFk8wjh/g7/
Sh2y18VujLWLtnryJkZObrFZ7S+2bVA7oqnKpHP/BQvTg2WbrSnInE/pux9LUuZl/eUhZpMg5gNj
+QB02jWcNBdVFwiJt9JR1BeKJOhjT245VEy/2lUu+g7/eMptImXv4qrLENh0YYHMv3BlAQB+MCdb
fS59yvL6HxT5I6NEZGtay6UoNASJtWKvfzmZPqOmWAKgIwVFNQa2q49Q4j3L7//Lrvf1gHLAJncC
plTmHoEMsiCWFRBRPXa9bh1l4CjJuzYHr0olMIqFn1nqu0yeIqRug8UhgSZ/GmphdwIGWi4qQI8j
vt6Vsst4trvTv2EOAQl3FtCUUcre3ry9AozOQlGKP9+I8WFUfdNLBFwO2Y+smgb7KJaKMsfORYPW
p4JdTRjArM9mLZBFPVj/Iaf2wqXYUDoWUVVEVWY+Bl+Q0McWLIwfYXy1ISqO/lKZE1ff/RVz6c7f
+Pd6Cemf6TmgLomUgWPNA2MXuYo5VgAEcQ94BqWaa65MjkN90dFjAvuUFwqNtHxhNzjPTl+Q8/oS
Y89ICcQXlrSTZsGvdsN6xLRCoKNMuZOJS5ThYQEuJeYRY2oimmV1TktcstAoswJok6w63HCT57Z0
ixxvv4zl1cXPmHscnkiDcg3BhHf2YCRoFf8A3DXEt6EXrRjK1JFFol365tPlCQRzcqPomPsh9N2o
Heg4q+zrC4MBGLTuhIi37awpazdE+HEyl8RwU47aBW7OHeOJkxHidSKsuY3cmaKK3qKJIGGCuTI5
ZaU8fLW2UAO2NqenpKdCYpynEHCSGYnVd+6sEY0DY0+kMRkyhsGVYcbfAn315WkooL9xzOKdnfXL
piAN0OKKNxae+cjmAEIkjbTB7ftaU1OrlbULETOVjrw4GOl7ZV+mzn6t3Fu7wAA+f4h65aXEzwGb
V7QVJXZi2AY6pY0Tz1J5IDHqCos/OeJrvLVvun1mdfvYEzyx6dW7dWxQOvMFphqvHFaDnddZAIXC
HBY4/N1s25/eaY8tgERQ5p7MSg5sivI6Kg/Dt1rCesj2qAc4kVXwJeLA/rvE65GzPumPv74bnshT
LPW2YCiqkhWHVxo1B/kUy01N4jWE1Pl6CFaiHfY8hPVjtX9BK3TyOGTRFsmtoKLDJlTDl+/xLWIa
zJ6zdqfvErEJDSUkQTdAjtcLSG9BITIRxToe+SUQQmL34rqnQzcpr6uwrM3d7tioYiPXeG1N5M91
HO7u5dxmK6gv87Dc3ThYIz4F2S3rCGDqGuldvruQiGqXIWX0BGxTAWoPc5qQaxLb5D5ANxMXUs/7
fQNdUUo6Apu/Zux1qTMSedWOTxfnMJNHJGxA8HoGVZaWurvVJMyTsNwr6UzoQa9HrNJ/d5eh5YdG
KI2WfAQ/GGljNj/EdZm+QcW5EPLBStYPbpYMgb798/ZDekx+NmCqRC8fRKIi+Rjswp0cjqjKdvRo
2nn8WrCa4Hu6sKH5+1jEZ/mjWuLezjdk89ec0/VkrbGheoOuyscu43hPDLGRJW2IzD+DcqtJVr1z
3BlpKmbOJJBmfQ7plZCuZZ/o2LyRt+j26rrfy+ZuwbkhUpvH+XOJoc65p5W9sC3HEGvZHJrxfWYJ
QlRl1zCQ4kDmUXye6+K8el0Ssp+NsXfktFBx3Ch6R8RHgGi4dMKmTt8lyzRRSrEDA3rODsyS8XpF
j3yUGlW1/UyWzA1AnQbonZXK6GfaqkO1C1cc2FhyzLwr1AB7WBA9XzTiRAl3P61zyKl88NB/LzeX
aCFVP6pTVfnXU8SWCgnEltAnGxs9GQFjblgPW9kxF7ksnVdHGfis7gHwxcqtYBS8mJeQutUJNZLk
AEsBcTmMsBnRKIHIhh0ru6ZwV1rWhoCX7W6FoYFxG14EDagtQFw5xAymckgEoC+hM+OYwEe6PVNk
LOtWf4+3d7ii7Z8n3LEuz93RI26ItMHuUOJ88fHiJrbGmntPL74MqWMacVD8AhgyWUqkgOSl1FSD
gGexC7YEcIlLGSl6maGLQrwfE7fWN+89rTkJaV2qTc6lq1aFZ/3JgrqKCDnwesduMP+/fib1wCBP
T/+AplBGpy2ni7cjNFmj901ytNny3DT+A/C+C8peuJTA9r2cxV2sIiii9mKN/gpT5M/9o6EeC4G7
Y5iAiR14JSmFGP5wPWSk6kynRVGMiOfdIdgBGkp7/s4M0TPsbaRuN4m9clSlWaqBlhtZsiF1Ov5z
EWc7xd6tYsDX6SPyD4EiEzCZPruxItQV0uRpAAne796Crl2JbXn8iCWSuiRhGwBcANDrukybavzJ
ptD1RT/ecPKy2f9Z4gCtIwgsAgbTgcuhLNmgtaM/zvoQT+3+sxfVR44TkhaSGPTXfPIgPS5WvMHm
62IO6Xj1Kzm63dw5TM9WnmyKFBH1XM0lYP2EEAaPHThmeZ5n9qgb+mY/9zkrUpZ7uqH2gCV2Kl2c
JWWuZ7dw5gdxHR9B+blUgxsa52jf+Izt/9PQlF18n6orugB9FviS0uhrKNAkeQwMGzUO1saFPoj7
0Du2GVrL0Ghqb91v2gCrbNFX2E3MHape0oxHIG+d29sv0cuA2tj10pRQIMlpObW5BAzOAS+ka6kS
pxJJRjg46xDZa3CKk5+/fLTCHc3lvzKtdKROoN7/U3dMelmqgJiJnTiIW4T4EwLduuJuv7nTZIz0
jN1EW8H1gmaU2xNHsXey0EGv5HrSmYF8Uu5MDcdM6g9FQEfLn7gq0Ht+6xTIwFDQ7vc6mMRQDzPo
k3CSMUcqXTl6RQAoLLDM8RAqhDtN1bsgjHXLKsvhT69SSzWploXF5zhhRnm4mJeGAQhlpyx/9nSP
4NLfIUccRTZY6Gv0A2hIne9qcYoh+e7/G1hW5ZA99CXIVMGhBjHkEhNw7N60bI8PW/7WvKdA/kAG
g55eLUR7lcSSI5DkXQ126pmwF3MSo0HcqDH9liSpnhk8BGv5eS4yGmhLLS7fwRD08gzS8Yn1ihT0
iFTO8mFJ+B3h75lg2czfUOAKcIPZmQ1weYzM5tgluEF2tYOUFm++skFM5pALbdX58L1Zcymqg4Fk
mVNckzk1evBclM3hgQka11dbPBCoK4mWJzn6lN4OJRnwM+JgSnIiAJiz3aoMP+G3PDfHJC9+pswN
70kmMY6u17Tx2y/V4mYQOAco4ueSIKkAiGAdhZ4W7U7wZPaG9jm1j8nRvn2wCmV2w0yjlEv9LJRD
8+j2geII8TaKvvRCM+6G3k5IGnUdo0NzP054IHVwDB5qLyZ7nenFnk5v4BnR74YyXeBU5AB/4eig
nkf7e+zUacYkauiUeI0qq4A65Mp6cL5XCWQ2fBZiaT+6vlu5uiINOtg18xqDQHaWuXJIGWKtp38L
GPNxn3DK5bKWAHCeVttIiF1xIOJ7QkFisCQJg1Brn+28Zw2xdx5smsXCS6/x1fjE13Rnt9+dd+q7
WHV48W2UX3RcgqjOohMAawYw4//gBvfoXL+gkhQcFH84ji/YexP9jxcJUW8vG0A/NS5rZTBM+aN3
cVmUba7vTV+uv0ktQPVn9Mm8u2J3DDPJKDuiEcQL7UwwHbOl9iSMoS15v0CPENABPl5mu0sdH4De
HqyO/BBj2XG138DUNT29Fh8wGr6yzfHBI2sQamhC/NPpyy2ZX9orthV8ioeZERI+avnlEmZ5F7yg
sclFA5csmnghQhMBE1lX/6Wp7I5WIjeV1IuiAFXQsjIeRIrn1ZCKBWjK5XTSTATt+Bsmexi7L6te
Vz1yd1QN5WByCxeTxYBi8aDwhQMCkUvrantOrhkhNIInHbbeU6YyyDFVg9poPOnso7SHmQwsvyJS
Opm5ICvRyIrLCQwH2wTd1JIBdT55H4+bp6Li52z8MNZAuhVrJQ2gimq87c+LECfOWZqQ6V2Nxbxm
mFRv4Agtj4wH7Zu9saVlGw3ebH9F+oZzE8WvEyWWyuA+IwyyK6ZaLK/8K2sduTmBbvbgajsj8Sgj
r7D5Kz8IMEzIMKVo2Wth4YQs/1Bh+XFfcz5c5g1QC97896VyBlopRG9etKM63hP4TzLK7dWWkrN6
3DY9FBbUfX+mely1llWCh5WE9aXXOSFoF0SawyI15d3x2sp26oiDUemHqUDPpJgRgnBlzTNjQgAj
7LawRMohfRxxNvqRSyQbsMsBRgv6HYq2TnIs/x9j6oe+MVL0FmHFDhtD2C9FfgFNnEAFK9poPN5H
7TeN9cZb3A+dt8brpErpReTvDmra1DgEsaFyRXiXun1+XF7gSDaKuPq43bQtQt+e1rqpJSmQ5vlZ
Gk2hHmuRQkJqEWu1re8GrKpG/Dmp8XSf0UGq0pmxiDT4NaSg4e0BOoCq8TxqvdwtsZrAXSQVamk1
G2HI1QQODz7Wq2Q9Mzlgtf6etoyXqmAq4JTOvE+apAO9+2ntnpwoKDAYkgSHbh6ra2quciZ/UXSX
LOf8hfZoyTPwvy9tqF3Zj02Gz0d62G9lRaP0Tkg5uNa1RoXnEXvhKYz1xKwAwnXuIiVPkA/MUaOc
uxYCRDFkzVL4N0bWEAGirxBcbwlx2sUCmVgm9n3EgHiS9LdvFwmSw8JXB/18q54figF34Z1PlR1U
u5dtchHzLYfe/Og5k4y25lIf9JFbdsNED42b7dNGpaFVHacZQ5W9gKYQW0VDeLdVuagnG5e6TKgp
TtvtFndul/XapQj82ifKttr2UGjf9Kf8Rkv63JXWQlKnKgcZSgg/ShCHdve+sjkQeNY8ftV1HntK
t3/ofEQH/zx5xfBjSd6GpTRgflLgv8P5Eu0xKA3ig6OpiTyNXwe5YJ7ocmb5SawtuMhHIdgZPZAu
kojgG4V8ApEuJ/xIU1yeeA0VYJvcWUddJadbQWqGkS6YwOs/Ru5zR3hnRIuq0dbvl5FhIqT8qiVb
vgRCOhxZFJXTQQsgnrWZzcg/F96/fkC/1oiCOIxw8ymiNLqBDEi7Ilxqf02Z+shXqIahVPwHtzL3
0iidkayWboO4INjIT4xl69cflttYsrO6wWjg+jBiPIDyvzM8dU5zlGjihfOa9NcdcukR3+G2ZEqc
qr8Pco238SK4Sq8l1yARQkuAbh+2RADS/VzyN8arvkr688Kt/6+XKZVhqAfTWzdmPD6NcKEonsvm
11M78mqC0TLzaP1aHw3U4cEPCnFDqnKjTOjRQ6og7f0T+p8q/UxTsS/SxdjvC6j2PdpSRjfeUneb
77c8ck7W0rRy0j2V22W9X/TVgKNR7Fxezxo6lvGgvWjr/I8MIIyIP8IKj6y7zZJ5qq38803vZWg5
Ej3I9Px/0M4dGcZB8UVAhfU3nznZ4ndKAUzAs+lqiZ+surfsQJBJyBhmqjvyTf4/p+CyK+jsgg4y
oGlmXXuye2btF+zZ6zerdv5toCw2V7jgCFlUP3RX/sM+bOzjMi/CF28cCeZ7vOUwmL9PfNZKozDF
DpxaU291ufy3kk/m2X+WXlmAAeY+zrMSfyA6IjQPyd2qF/DJ8sV9XnaRY1fRomirb1eNLXUTBGeJ
zeLp4/lSZU6eqtTVOnAEKuZPIEnm7cMkRk9bq4Lt1CTcPdTHuZVO1V9JYMZxt+hfiDZf1KH4yyx9
TU/s+M3fei77RFGGxyjWKxckGNIAIedvoadywD29axYaj0Ss2SWeQE1tBS4ovACTJwo7l9LrTG/u
GEzOSntqsEYe/R6Lq6rlYB25OcMe0k9bJRTKgJp9SGyfZoUo9HXSWv4PeQcPY5mNdbqlhF4KEgAd
xzh7Jif1b/EBRJCDqi3iXHqUJ2mvRu9dfKA7b01cEP5oMrBUIrzJt9rRDW46D5yjzRkQVV2CTOeC
Ug6gP9zYY+WliiCkgvBICHdJiwmUKAlQ5leSbDe6Nakgm1CwnpMl4qgrsQQsDswd45byF+WZWrRk
xjPnPSvhdz+3Q6UIytlhpzvyuwYOjQtbK7Hc+no+/y+OemaT24QLlSEpeF87Tp+OCKWRIT66nOSB
SJFmlWtFwu3kfAECQnDHg7NRGSuKSCjKIMTKl1nvgZXFKDeEJj7rXpMJ3bifY8pidspztb+oQFZg
BcaniKUBE0cYFchgC3++ZO4iln+dPyGv8DE/vsl+sL2EcqOIJhinFp0jU7bITgM/7ePBiYcfPiFj
FWknp5i60usCl4mlj1LmWETtSHhri0GCyKwuk+xq+yeI1IAxub6ALlcJ05bI84nqelUKVp1Xrm/G
EgEcqfBqu6xgO3VmgtUx6Tu8UTcrI1BtGUBvGLZ6G2gVx5JSXIa7okBwt30ZZZX+oNRVeuWkaZUj
75BIrPnVPMimBTYHYalj+fbMEEQbOq3c2Vef00JX62vR/1zD2eIjOVUY+50qeyJc2hACZSzGEzFy
xnJGPSk0ATC9USfJr5Lsi/p5fSvNs5J5yNdR1RmTtm5aXwHvBnE3ojnMe7jZFT5e4mor0vz1HUdY
3bcGI8fj+6403NX6zlRvqHyy7vaJ14DTaRJbI8HdvLq97lrXR12tdTYbCBL7jgf9AWgO04aEksel
KTg+iB10w+3daCdzoqkuTJ5KWummvEarhdG8nnVKUOoae5YN8v32sjBdVafd3FRTT1jX/NEriphE
ianbFN1ypOFAgn8RZFz7m04ll31XtSvUt7gYXlRNkAT3/628XWYAcH93ca9wBbU1G6YXlj8uPnpk
iJZcpYQJhfGuSi6/Je4BLpAmaazP7UtVdzqZv8oS0Eyp8UdaaJLCOFG/EqXZbF6Ky1rg0wdql+D3
JbIOuLBn9tn1hhg3YzXMhPtve5vmNRVgYIHrjxIg4qdI2hiIOUyxw2WimjMubTSra2f8hY76AcQ2
CihPG3rcdR2GoQ1rLp5saFtJpQ6NkB7LcIxTzJWHwt9dz4NxmIiNRNMc+TqwWvfbc66a8cNYfHZ+
X9WDBcaYPWqTcnx7eDPrWLSnXyP9t66lLfoXK2obgey2vv8kqZgV4td+wdKmsoLXYxAD28GGwArS
s+2+ENRcB7UtlYZKRhGqMtY87oLXXdZYEHs/hkmwL/KZjYd5omRSeewWiMgY/+75AwktNR2qcAvs
BC3/NTwDR2irQmc6Nds7uV3GWQoLAYEs79FED2oqIzqbOvJuZIA0iD7lNcsOP0NtSRY3Gxd6d10I
p5asnOUJe+5OLyiWw6VbNDD2kgxcDSV7/HHYqanA8jitEBCC5+h+RpPD5Wz/dkuEwGzPzdprUSY3
ULOqyiPNZ9Vfv3FJAFsio9ixq7Ko+G/znAyRwe0l+virqxUs+l/jaUJ7do/szQSfNqduQutUnjIQ
n6Ud4W9OT5ejTIMB9RYu6tgLSBvEU5exrb9RUOuNiEWe4VNRkiG5TvMwURIaWU+AWlVm66ic6bj9
leVUG+8ECfhLKXMMzP6ulNH6SBF5yPFW1ypWxcRfQTSUZWDTaojNi7gxhFGgpxhG/ExQeSFH585L
b+J07i8+qi6SyR1ch/+Mke4Uts4Ef1IbcMP8lybP7+4rQzVryuoXDDKjnDuc2bhvKLic/VBkQLKD
3/cbWYj5YB3ah+hwyivDo6myAaQQK8xZAJBXDOn4KoWq2oVvwQlphcXHuM5f7y0gnu+jScUKSmMf
bsR6OPEb9aJ1xGqhKT1c/miQBHq/IMu/4A/ug6+9Or85//N0QV7XjW58oXoYrVeC0KYNfJw1nl43
Ch9evmWmHVFOW99fL6SO/iyKzm7MpN17c8wN8IMT3Fv/9cByUV83IjCIS9x021A+MYTSYClg1r9O
B6m7iGQy3QLl+441m2nUask8FW1UVSwmd6d8rN9BfA+AGzs0hqUa2bg1fDD39pdQWvrmrE0N+nQb
Zl826OGIEJdSIpc96AN1KVNOlOKAN3+p+prZQPR5TvUZRg3FDda7PtNCkdqt7rhJPtOJpjVnvCke
jsRewklXyQisdkX3wsDOd5T0UCDyIroo7FzQ7cwW65G4Zn4MS0bATrC/TcKGMRzTLzIzC6tCj59F
9S6v0b2BGgVDaqDzCujh5+Vgp3MHy8GtKJuEknbxYaZYjnRsQLENAKdw2cNkXEBxtt1fSmnKoudA
xetG0BA24NdWXiFVT3QoCjkzjmV5j+NgQrS6HtLvKtiELvEO7ohT1YdPXiOhnhpwVLGpaZihdNLc
YaMmAZfWhKMcJYwrCvbddYkex6iYndsSaHfNdPFvwpzS/by2Yly6Gz/UoyOrOaddl1+G0OVxaeag
wGVmdyD1qgfz2plS+U9jWfHpPzrN/Nyxm9Ax6m9y2lWEXMUSn1c/I8QaKxzOiIKf16l39ycSmj5A
S4AwSlqY4hui9OXtXdm7iPdaVRNP0WZWk0GV727R5Xy/7ZB5WY6qwMEmNwpIoDaGnhvtvOSmUwHV
5fWRd0B2xAvF4RJxNU8z/Z2hwOvLoo0z1DZ2b/91oBAjs86oX/5HvHajNiOUkUiYiLng05PRDCqk
S+I6gVZkFlcLskRJ8U8MvTbwlCNCy1U833RJF66Im7RSSCH3zshT9jZnPlKAO8W79iZanSXvZECX
58NoTAcS7Ibu/STvrlAuxUJTZAhik/mIfDlJbsipysI6qxHKhTpH1qU2eVgSMj8xm7OL91VEY6Ft
RnYwl9TVnzwmasaMDSe23ZLZ39D/r6lItx21Qg0pnI5WtejySoX2pfCDIGHXZJF6KGMy9x3Itu5l
T1taatqOnr9mVhezQEEF9O6oeDWnujH0/Q+h2Whad8MFirmGJL2ib1knnOPZD4fxBoakkTUlpeL9
0mlLnhQ8aUpzmsGE48Vp5BBTVO3KVD3mc5LIl4xl8FdDbJdH6qfdb84CD+i4iokH8Zq+sY8tSNjR
P2RUx6eI94ZnIJtXX4POXiti84ogT16Iw+SzfG6XNk+sd774Ae9cWpp9r/+0bkXwplslEPIGYNaL
2PcwxS7RCJE35ZX5aWHsV60UD/wIew5FucmpS/s4pTHsf6Au7VSrSUwrUDfThKBH7bUEdl4ZO8Zd
vxndRzqO+75azFRKB8ixdB1UOoF0LkhudW9Id7ujLrBRqhk/7EFh5134q+H6ykDYZoSVRcaNc5eY
buNGiuvBJWIfgH7lnSP/hhW0MBeA3Giq1tEGt/Ea46Hx8qXxXi5z3wcDWy7qTkpgjDICzuTgOsS0
wSVsbpzliMc3yychCE68QHyC678DydeFFdgr5sy0y3DnYEOSwfYL0AwWMmEXChYS6GdVl86a+UVa
L2C/5wj8RpSQeFnZZj2mfUE/Y6oyq4mfYfyIBD36/u78VNfqKQHfeczZoXFDpQB1CFRbd7R5CZAC
C1b9I9ZOLvdkaiwlHqGn2sAtAxc0NJ2vNXk5nomaI82Rub6wB9tUQG8ZPEH9W0D6F2Ht6k5jzl/C
G6KyNE+kzIb8pw4AVQiIN8YtnsW19pvPF3Na6Z6xgLZtsnXfIr5/Eye6F1EkisghL3UzOcXtUedl
R4Qh2oxql7Vs//9e8yS7bm58nU5y5tgBqGBow+7G8FSHkbfMpu9rweIXHKpQXIFyqah3YyLwk0EJ
hqLkupsgeFosrOz/eVkkT4m0Pc8vDbO0YVeDIwrW0GbVr2NW+h10OENIhPPFMYA4Z02ufdztpuLg
8eSbn9AXssQsOw3VZyvwB18wcuTEDbyec3mbOTiQvM3Td7nQ6HaqII7CuFD3/D6wvKJgOs6Er2rx
BDBAvfrVeepvEyZNHD1sXhmvpMulk8M04YX24b6/XIjI/mhdJtmvpJVAiHK3VUVLyeCtvleoNON1
KHLmE0Twl4z4ySvh0zfXjL59Vt/D5ZovF01SpbGeoLx8fzCH+6AvbaJ5WxOeA6qHWu9HE/eW0b7g
1nE6JFrOkcyHClWMyfqEq3i2Z4XPg7/db8QErJq8c6U+2jwEFNGfquGYuQTz7bChFyFP1ZmTRTVe
PPeBhKCUbXtl9iCDk6NWfkIQY78GKHfmnh2tOGKpwwBqD8xwXmDLMDZ/DADPqZGNBhzurtTUgf3+
HxPV710st4axyznd7YxK9PJnkCCE1TychjSsRzElIDnhEdJBofEOxNIeRwQG8inUS2hF5nZWQF3f
XReBr2HF7CjL7WELUVjDhg32kB7HOguAP8lupsfnF6ATjxEMBi0RNKlHVPtK/RaPFvasgOlt4Cou
FzbzOFFvnmyz/1s75ufg23T0PLs7Jl7236OJsdM5MOY2wWjZ9n6v4ynWL1jsRC9OA6ABoBDubPcy
b5e2VM9IHIGWaZm2eoJiqF1TM6iy9HmuxpFjqJGrPF6kdA+9/uZqs1oO4lM/oAiLnwgWwd2/Hccj
MjGp0ZrJ+hjARgqm+OjxMjUXkc7NJQj7MZq5rdVBb2VuwoWfcaqIin1VKxogUu2aCFRUesI9hHh9
0P3IzSjxDsIymnKW5Yc5rb5+aN4pUeCbPD1Vyw3tfQo/oAOEpkNGnFrOr+PTLYErHh56+I0v2vmV
Lnk+n1LxHsd7h4wZKPirQuc1ZvUBV2wkOUM7ZMEAfk0Jh5mGYIgpjCVWrpSriHOh9GUfMCxHSG67
xwG+zXpmZc1272nXnHrNTZtC/PSDWuYG2tYLrBCk4Eqxt/g2Z+TqwcLw9EmGHzX8FHlHvi2TcpxJ
2CR3o74o5dDcnnfKGBbVgPT8+TjYy74xst40r7F3PbJ+iuBzsCiNb/+Js1H9NNswcg1Yxo8h/3qE
fmP01WhYoZSI1Stj/tPS17eGH/+z7S0YS6LEo67eMnwGRS7OPM2v6TBE0TIIVLHo2s2xPEXXwsvU
KIJ/4ZXXhikE0VbBsPy9v/zgKiiSVOTSgsMhY9+yN1d/9iCqun7P6xwqWh0LaomYrnXkehtqwdbo
FCSwbDBNmFzJQX+QEN7q2lFMO7GQQupCXcwyguU9YjgTA/236iYqsD9ZqNYp9hby727etGrvx37Y
WxUIsM2ZQ6qgU1zziwDiKq3VjnYjGw8gCis5VwYfFY71ckoXXEPeCRRXnGRbU5cp92lxLfQ1YDLR
8JY+RjPDK22wBknNFNUt8NgFIvsdfYBp6e8Gu9h52wf/rTcL2n7QNwkvov/BkIFOQAu1JYTK+IOT
WrHB1uDRdMdE5UCMEUD5qf5tUrISIoUJgET8aozt57oSHq53sTFvP9T7uBYfRtWoKOF8KF3KvL9x
1BhN442YwaMH5x5RNNTlgCTW9JYUNsnU8pTOEl0xP/GpAng3HYGLi0kBUuVueTkuPdKs5mQDb+wA
B24UpmDG1R/xpr8yvOlubNAaI546FHj3aDQYzv4MgXMsZn7aw6aCFhJMlERZAynZN9Yl+ycfKtFH
QqbHRY/Q+jL2rJFTLkbvYNWIpySX26MmAdseMhfA10rNCpK+2QzMlAUdKinNi17LthBYtCd8KuDN
dxRvxc8AWMHs8RoPFJXvAmeJho4NveG+cn/PlAtGm6XSrZto2h0B7+CP88gcYCr6iQ4VzKwNvgje
bIF037eX0Qc2czU0qXPfjIPno4f4wsTTiiJmkBdHpozT/190HYc1Nv+C5/eW5a0j6EnB5+JN2JSY
+VPXxHHC4mAZ59WSZeU/210aTv/vIXCqBJHkhgIHBByDaTacHlyEsxk2sVPoYru4wFa39ut7JavM
vx6qbz9/qn2mxPh7AbeaK+YxAhUdvmkXxit5OiA6/p+wvTwPtMJ3uD+4Vd8TpyEES676qmaYFFZt
vQiCxMn4Y3o0InQNkuw6TupsrCxrmdfmBgxKYvzVYVWjFojUvah+6kqiQqphpAP/EPwzrGWYfdB2
XASFYDY7T2Q8PfmQ4eMNs2qnVcRLysLTrmzjx9r947LfXcjHIuK+x5w+O0DwXA1Jkeo5Qr5c90KI
z2aKGyqqtG9XVt+gZt2Lnun7CQzVH/Ncx9egCO3yAI4S1NUkFFPcnXe/8sPgQFaQS0ddmEMkAtmo
9mIPbsxTpB38I9VjGwQSCjOnzKme0dXURMfczALwrIW2B4qGzhBE3fuV1l0cnNTcCcMzW5rNr+4i
kpjqoW0u8fidUpSI0otNl7SMtfyiQpfQ9Jed5s8KNkT/gs0RMjG5KlcUDpGifTphb4Vo+pVEMcuy
7GnFwdV8Fvu9zrPzuXpzOd7cvjb9ot1x6oUcBOVCziPZduEDuVmd8gVz7qqRFzy/LnnaZYJ/vwVb
gKdqder6M/qFjR33f9lNIg9N7iHOcJotJvEwsFJBV6U80WDzhcA5n7UBhalEX52hGJKqFz9+/NCH
cj7eAXHIn95TJiEMf8LlnoxAcC9UFDH3LgCoHC7lDT255pbfoO2F5y4NGDRY5vR30xHiw+CaHs3g
vpgWY0JRYzq3S+5JDIWr6tUAMKtylBrSzNeaa6K0gmT45tVKH8v9OAiltrgRI1wXHm8nHLeX+eZT
6yIkA4+Z4Ibq5AwlxP19eej1iPkAWRXZi6SZF3tzZcMynujIZVdif9CbfXlcxS1TY/CHrIzFsvHo
gGlOBh1z+FQ9NzYk1ecSp5VUs7U6Zme7qxnhlaKZURQEbITcbL82vkCZe5CdHwWGEfEYJAfmV/Uw
5rpocWy0bxX4cUfjP3D/wk7WYXxlFiT6VomUaxhEY7fJUBZ2Pa3dmrxcx8yegcJE73wOjJinNX3a
13/7hP9GRPy7NvZFpnlzCYdSos6lhjdrrFcPgrZYhEIJKqT7cUaETcjVyTH/2KGFZlTXed5Wu/Qf
6JDU5I7H08bpkuEGfqOv3BtqEXqvMc4U5NMWnPrQi7L/CZ0vJyvnaU2CsVV/nIGxXFD2JW9pXYi4
sunOZTwLFkrT6LTP1HfyFCsrLPsGZTUnZqsrPa/OAVwiuar03pw4dL3AbVrs/UwkPldgqhiEN2sf
8u73O6J05TQ4s7qWcRuvVlUBpZ/bm9RVVNuO61heukNgjt8lR1na4vHLSJPkZg8yMkq3l91DWLtl
yZb38gdL6UxzhMpA9B3WrGmETXuE128Syd8GHzfci2BF/zLtYrXfqUyb7YLQIy/fsShU+ixvpErz
aofAhFfC+FTCMEGq+rOkiBZFWk9yCTsgfIUgu+RbXuNWvuIuCCRex8WwWXg7fY1/C1vHNJz44Ylg
0eUgZ1PbHbUWasODkHjH/izBlA+M/whoG6zW+S7hVTaOc0ZS/GassrwEVKWHgi5tNAVmMSljozyx
e3ZFjrNbegf5mqzrv7xIBtG7CTazYOSLJbzIG062fGEaSxv1i6y0g1EQWl7/Gbo+fEEPrd1ErE6M
n4R+4ZxbQXB4+mUOsbiW4K/+0kgB3pm/UwHaWKTYngNkOzOeT3Qos4XbWSMQEkWOu7Kx1hKBXDe5
MpEDaO1w2qj7ZT5aRXdfIzPzHVZLc7R5zLctMDQzFMw90KxVC+ipwofg+sYX+0rovmbQe41vwwau
3nSRx03oevvPrso0tva4YE7oq28pE+covENCGyMGstrvF+swHi/CbklAkAI0JTTT1YecuHe7k3wq
u4lqLb/Xe/Ea7tRufGFjuQTZEQg06x8FOfLI08ebGuc49LuTMX+3R0y+5cHYrWkG7hfmW5ytho5D
8Kicg9Z4kD3L6ygMxcGkZpE9XoUzvuOifgPorD06JVsfpzsEmHHjOIWJMErVloVCxK7CkSXBRdUQ
yp5oEVDrLh/xUk8dk+igAB1Qt+a8cxcRRVg5CmI4+Pguqa5JUk6/JpD3fxDYADYXkLVCD2fZnTAh
cB10Dz/DdVT0xazUE6iKJW5jbSYdjAVJSPDRIXEWxWzRKxSuOUcpV33O8Lu0aB9sc3aTUPzMJfXW
50EHsAtykUJjy0Q0h2fMtXlwe+kb62IgynveIVkgVWVF/C1wnOw6zZF0IbR0rrKlG8LMj9dqggik
TpFjsa7Ebs/jYBd+VjvlNhr4zsFodD1P+LvaPHVWaQrjq4uU6dO8fG0vgrt5bsKaMBm5F49ZeB7f
5/pyA1DIov+ahorDmkMtx2GUSRLcOVENQJi6NXWnUfe4/aO/UnIt/Xj6qw9i+xG52FQQGJH/h3u2
WUvisRuV7B03ZzGRMv/XOkZi9+mGbgyDQLsFWjgLWboLiHke4+P0Lx+ovSH8akRomTbqqaMp6vnm
+sBYe3qUfYI2Hx/WArX0Lvqh41jAEUj9958t6xD9VUal8IE2UP2KmlaQ2AjwLPem7Y+OEDKnoI/t
hKerob+QY1FefEKDAC8dlzfQAJpcKdSLgj9avdqZXAEXd50cXCRIsU/c1+IcVXslh7kH5Lh556dt
K8ML1fGQY7Td8mH5uwX2tAmJ9Al+4Ri3sLbTA1DQvuCjnhvZYw5F6Qz2lqgUh68oD3n28JEZFOmv
dakyya4dju40RhOJaii8W/SACcxbWzkEOjZLa8m/VcIyjuZWZtR7e2SgbMps9vzUHwL1b3Wbl2gu
cpE5df0ZrG74+KkAoaZKYLtwgHJ0PO4bmH2h6dFb0+y8HnBiU8TEfQpWhwPTd3gPvlUKAbDmTweL
F6ZDiN9q+qQeHTtqnt6KdrBE4jdV5xLdIoc3suI7P1N7ZnYb1o+s7rI5esEbTvGPlY1z0h6X5VjU
ADM78wg7kRzKgMTYyiOY4nrX/8dIorBSGe+s9Hr1lgLILIxtlTO+Kh6k6mcW0EX/2RycDTbuWR9E
ZRb/INAPpxbsBb0wzunK9A6Jm5U7phFOjcoZAWxo0U01Yn5E6lRDlG5s6I+m87aHDCTD7xGyVR6z
Pbfdh07oyfayjm2+hMSw/R2VAOo5tMIhCImmgg8RnRxT9b+/W/IYT4JlJwTK0u4HqCSmdjKxhbAD
a2T8kK7lHdpitBmZnKmSX3Ryzezf1AhNNcvRbpRoMH5ASzg9jsQdb6IYxQnUdKAulki5mHLfqqNl
KXQ/w/X+a0F8HzgGYdlyJAA7P0WsvLwr5jreFWD+2ULGTUst1IFszFuVB07WQ7zma60vOPUS/hh4
/r2ilvfwTz/s5NlJilfJXZgVf69iQC/p/l8/VnERI8fOb8fyfogjQTZlNqN57nl6UKs9Zsepd5A2
r78BLgh3wSrwBHFaRaX4QcLclTq/l3OuDz5PBchiAlDU07HGugQ0RXwYiMeYMPgGKekSxkQRTCKu
3E84hS3ISvY+oT8nkiK+cl5u59/v64MKY1yEMkDF2fWCJKKgOe9w0SgHfDGL/fxR8MOBOWtpAZ+N
TVW7BpThBYv9CyxreTAMoC9oCls1fKOigU3Hpr5rdBSXmMC4xEzYq+eSUxF5cjDu14o50yGTxLLI
USrgzkxTkUmQ7ScaiqVgR4ZK6X7rZkMZymIw/InFMoReikQK6NYv5J4ouFhtuW82Gl00N0HeRX3r
C3mtvzoOyWlOLmnvjPoXXM73qhDlx9cy2SX/JhFcFejD/y3M76tRxz6A5XDSvX65HndwBypW+nv1
zjU0FrlkICdjl84XN+wBiuqelr8ncam0pj4eQOzOyisNvdk/OeAGURHpbilIRzARc4NiocXTVuyG
MSBsZgrcg7K6QFGHG1dRb/cVSiWeBr/DK500280qupQUwVg+0UVtUYnqo6KbWPhiJLaZYVhmnm/B
VEcn7xwqQqzTKIKFkxsfoRV3AZRkoUJXohT2GLIWeum/tfpQIjsWVxQ0QUUD4Zu7VnpVwGehiZw7
M1ucuaHmLCvzqoPUx1m2xy6Loyq2I61pneRs3LyOpMLcm8q6dPtTJLygh4hukk3JSKuOpjpoBT9O
v2PCXFXq8iKPyX7Et9Y3EFflYDy5G3qkcVjRFFrLEyFVXtLakzJoIMZx9/Ztx31n40k3KpUuLjva
dk936uopM7URKxxkjJ5oF8qNnmnIfAfR6TNB/q0kOwsT0WQ32keoedV6rsJN5pt/DUZUohn3Prsl
tbH4CfHH352lwd9zwfSsXL1lAU7subkt0F7JVcD1vl7+dw7rxoNUi90rd590pErGYlnbROj4B7zR
84zookXrvjY0yuu7k1hZ1J3m2Zd8W9/brJnJRtXX0RB3um3VteaI1OtVxpCm2MfLX4RfW8DIQ/xT
vG0FyzU+WE0g456+ZblHpzNIH+uyNKwcIChUYwVn137f0MkXKC30L+oM70gXkgvx6iK0LOhlZJ0S
WahtuOaUaBSPL5vxX9wyh+KkyYhU+GsASKKW6XPj4exFMs1S6XQ27hypml8nwkEYLsCW0NZziR6j
BhbLKUWP8gUW0V91roKayR5WOuhrifK1boBcmjJntmFuUx+Rx0z0nLZNkg+d62v6LM+92lGmjcYy
GxuKa46Vsqa8spVv4F7T1ZBr0EkhIB67wD57EF5vJoZD8rSQAT2sjDL/bFau+yuQRPz+oFve7ZVB
KB6mQWmkO+f1DMc0zyFBYkmqAhc3gYjiFzLebK7wWtM1kfphnIXa0mxTuKiTy/0QDN4ND3jMv4Hy
yGIU70BTSNTTfAhnUs0uTZPn/OV3W/hkCRCe/sXpC+k49uYbEbdShN8aQsV1O2nKnTUS4u23/3uZ
MgURnQ9x3Xez7bKUaeplUTn9SYADYblOFHpU0gOV0wX2meN2xoT2jhx735zP+kAYbRxb7WHZ5PQj
8IdsAA8o6N41H3lX3f97dspnS9qAfASFnmcXvaIVS8wWFWQ8nbw/jIAEZM0V7gd/l21x0VAmMwhT
0bEyKpVJQUAzwBpFoENwInH7TDz3G+9PQHoCw36ItyeE7X8zN15qj2vZvPR+/UhNlsk/VJyL/CuU
sydykIPWsu7A1ImDF2GQNocxPVqXumtL+BaS9IFQTCPoWYXR20hhNeVNnd2e8iMrOduqmI3it0bF
nqcWgMevUfT4UFK8sdJFTE30HOcARW4UdeNUuVQCSJDlbSjnuVaLCjT4kZQ+QzElEwIJ6DmsiYFX
g/uGg8YglE5F6UbbEjJQbmZ21jQi//PVdhOToNnPCyPyPz5XmgdSsENPBc5HrswA2iS0A5/G5ZO7
di9g1Y9S78osTxyukDtyAhn+WfW558h4RjIYqZ4BCC5QfsgJ6jwed+i7dyn5tYtgdJwlHROQo6BW
lUuUBupH0PptuzxYriX4kUY6/NreGKTPDX/ufMt0I82DCzbA8KDbE/qo6l6uvntLahOyMoptt9np
5aGG/rrMHACEUY1t/ksWySYIFuNmTmwKkDFnPuQlU1JEohpIWr7C32/yeKQJTLRJNXZGomHKjGeI
/aF+Ynrkk2D9RHqpVS5Gf9hCIXA9a/apHfAr34fFrYUd6sCd5Zg0PT5ZiUB67aCcdfPgl8B2Zgpy
waeHlDlLWv2fqtav5NkAIDX8ra3DBYzZQBlZtP3yBdIAlZfTiugqRvuQppQ5SIxn9Iv4AZK5laAt
T5GmZWy1Ozp8lI+50hy/PrnYYJ1ly+p6G/wLvoYtc6wfyC9p15cb5L8SCdF4J0R/X7/eZRuRKlJv
AldmRpbu6R/4WjbL4UNXtyoSkZcJFDrzEezd0w+DCtbakQ6RCE0w39+JGvdxDcMKf+pDPlXq8kjs
CALw2emPN9aKi//oxzIPXKEdalGFUx3cc7rrvi6ngyljLzoH5x1pkaoWvdAHGUylRJCPOyZ3OazV
9/bRdpMow0ozYSYCe8EJfBUkYao/oBSkDI3ZbkDUdGDXGJscYNPYr0YDkqaw4KX2DoOw/M+OQT86
yfyJNLLLoiHYQQTPYNlcVTcnwjrG2BTLGsPz9yRFIUXAORuACLPUkp87mf4ogfrnq+MT3R7av5/R
33By1BMb40xGTYZ3a27hSSd3ysHSrtwa4SiJrGwybf6WM+2iNSBs6lADgONCJGp3Ddm0+6bSNvXr
dnPXPq8AdnE/LeJS2W2oN/NAet/970ZaYBVFCrg9JaifPUwp/BqIwoBYfy23lhEqPIIs9ArUQMBC
0AojmevavUqBEhw1QY6BjnYH+0ep+AUvZDALYUEGTZNOuVzH5Z+5Z/g0R0GtMkXsxCueEcmV8Nfd
9SgoZZ9O+yhxZDjQK4xZIJQhabINblmWKnC7bcIC7whBJAtfa/rfM2h/6hEMeLnI1tuwYypYZ+Xk
I48F8ibVUIhLyF+U2le+n6xHrY/yR7+XoR8E+HS18DE3c/BEUqA7Hcq6RUTqRIGLaUT2MmPDWIRo
rVzKPIUPcbngy6mk7DfAmcGrtfmidrOzFBuUnSP+ufdaSsn3nXOPDx37Q5qeMEeWHvbEGWpnMqUq
d21zvPlfIUYMfrQ8Bcb0r9Fznwd87w7oD1VNT8GB8toUgwpOsKTMsZdyh2Ug9Qg5BCcy/9vMePrL
het+5V8qpqI0wpoRUBHZwsWhSTMO7bWQpmbixHV4rloRomErg84pMU/yYoMuH8R14w6YuWJjUs7h
DPzCeyo83Dnbm2YWUi5T7jk8IEyvBnfMFQH9mAFWAzsdWuyQ+GzwDDH6y3KlSa68DxXdTOjGs5e0
y8GLz91BtrdLPc+xz7jt4kjTUyWAf90KblSnl/Cc845mje+Fuan7oineUEr/oVKrrQ3+uIV7NkOQ
0+18s0NrDHN5QdEByZS3U0vS0+j5ktYLaero6TIrpVoowf87gewhJZX1RxZ8YxngXyY7ZxkOchXf
fS5NeaGiDewtvUGiw8FyCR43lx/b4NCTJPXsVTfHMnbnJmjaki+CrUhdgCGbA5W5Y+EvpXg+owgF
M2s6j1T+OzgR+Wk1EhNudbkSeqdli0upWris0dGnAdBMm/INWEO8zga+x1RoQSmUvhLcUfXk6VYe
0hEOLyEd1oanwAA7AyalHXF6YpYk1OnDLbGbtTbahpsYXbGoTnZPCVXksSrBeivVE912TWCx8CA+
4Mp50xRYh5+hVTFyPl3RO3tYGl7s7oH7YAF8Bc9qR4fkGvapq8ZTBqHeB8KzQ0rSzfqGVMA1iZ7R
fFaC72/IbjUWDGvX/LEX12sxyUvN0VFx46jY+iSy1ufd/LwKjwXx53ljB/w0N74szcyMo196PGN3
7AdBUTZiYgUCB2vOZV0T/uu7oTwSISyIHhpQbbgxByrga8R3TGrCGj6NARFyZyRGF/6E2yEE6P6V
Q5a8MHgRoZRfjBr0jnP/y5XNmBMZp6ko4BDpW2oXoIpN437325XpdVvlhPze02RdLSowMSJE1Nkk
cKSH2g1fXM9nGWbtgMu4oM/AQczggSla7o4WkkYnlrL2wT4bKT5bDNzbxQi+VZZQbrr4vf8SKYw+
WQQwGlfjwYD0aI+QnCqek3dGjy6MDHK5VqruK4PCuGoq0CCLysbik93jR8B14GMMfyxvjiDc7DGV
UfGZBxVddFCwaPT2if8BxcK7e66vvF7fYA3NsiBrtmoGOS7hNOfuDQQ+Ub8hYlUgykpOAi2iVdoX
La8kcANQn8yfBtqB+xU+vk3/uxAfpzlscyf/UNXFrptbZg+Ztd6hlCe7iGsDpdb+F8KHodwkaD4u
5MEzhHEI91XZTRmnAeIaEjUk0SCkDJRhpgD+QvLFGGwksmeiJTcLadJYML+DX6sVDlJVoOn0n5Cy
/A65TWeLz4wCIQlmef2+sW6VcffP4IMB1P1X2NZAsrQjXu/R7aJ1PACMZQwueZabUJYBe19h7xPw
rzjoxH8tt2Zp/+pRgFOZoWpMFHP1wvpCQnTSh+gH550slfCoXcJDhX5TkcuZ2ELteQdvOyRbcrgJ
4LLWixr2jLf5ioqJ7vspquqrnCW0ynMs+pTAF9RkDvqUAqeHlI11mhrSr0DeqQdW6EpGsUYMFYrm
e90OkXVwYRn2kK3hh6Ne6s0B2Es3UZeC5ihONqNvJv4swcQUwsC4IV4WowmlipzEp+t/nc6JGwvV
PFEVF82L4hw3x1fWVbjepkpOgimBBHUvsiILXMIhdsvBuTeFP0VFG5mhb/O6N0f9NcSPXlRT4Oi5
N9H3D5nq4kYUhwEeaqBK+MGn+H7at3i9ASRnjizTKkOlFW0gfeztC07jTRN3ODUgcamZ9u40Px/5
cBCZpIyGhaWKifJLSW2DvsLnzf3nT+qIqjNVfSkj5DeT0e6qlrQJgYRiw1eBoJVtabocpkiHFHa5
8E6MEMgjZwiCRv0iSxn+pS9OUj/IKhcnThlvd7GfY3aNeQp66pOjnA/nndsnci1E45MTL8PEzmgR
IgWv9hpnuN8rGF/lD4OHtDgDup4Wv1d7aOOAUBrQ5EqxihLKVNbVkAEqy8jvj14+RVPnp2kFy9aK
Dxa5EctijGKUzbFytWCXSav9eMoFtGJitqEWCVDAGzp5jRrJKqwZIWMdrHm+GIZsw2nNI7XguSYe
I4Oo7iErGyJEK3AlRJ7L4sRgGXBg0H3PIqAChthSv5+5+aDoBrCm/LJjEdyvDdn7YkXjL7Kim/VW
ZbC+V0F+hZrs11/YtHDSUBd/z9TLZuqXdGHF4sQklJOKR1FDvA/ijEuQNFtI247krayfOIcOMXen
HbLgd1fhjlUJCJ8PHba1JAd+vR4X+WSbzHlUn3e16xnsmjO/jUuPdSNzvh5SSOpLVa6JMf4smLAB
8EfbZ4cX27OPF4ym7PfJLvZI18ssRCyeJWgC2mEUpAKaqDbI87DzSSOFnbZHU8ooYssIOkdXgF36
21DnA/VMAGc+5DGk1V32kiORG3Kz7r7bh357+hmSqPlMUjuzGJC/pvDAeDVlSCZsfrhoxbquwJ9l
Z8r7GC1/AcDS7vwstAx3Cu/Z1KVrcNu74fIrCtDnKZUnzE9yIKYwRKe2nsx4yyi0sghviZ8kokgK
jZCBMoXKzYmXYdB3OspICjq0j3x8WJidKCmBRuj+qQUCRjat2oA+9vTKpCY5gREF8yCAMe9Uf7QU
8s9TIwlUEDRp7+NuG1kPBayJGGivP3MdbZdyrWBN2+n/KQuX+4RfgPISSHshXSXHiX5D0TjBRaPx
XWIVPiQB+zoc/YfwlDjZsOzUbJyfRAmX7xEMG4TjSF2TEvdvIFbYqrqtjh60ovjlxWfZKDvUK4ln
5Sr7igH8ORSglbZE80quTaw9+h6ZX2yoRhE7ivI4sQFrc3id63yB6mRS0yjIvbbbfEIxJ3JkjSro
bdaZYfOZIPFbbv37AuV3NVL2P0NcL3qzrMQSA4kBOQv1YIsx7GGOmYgalRsDjIGgmioIKvyQ+IhG
3bd9MwEFzn+7P9NQKXO6Cetqq2RJYeKs46j5KW7bn9hMBcB4+lXWSW0JJO57IYpmk7qSF4G3cshp
KDaSQdIOnAv5/bwPuGeL8DkUBTzSHcqwPEMMT5mAu8vAmnV18WR2JWRcaq+bT5maqmXK6ENVB7bp
tc248NuA/cWXs3B78bt+6rviXdR4JsT3707cK/oZ053Q4enG32ope/5j0ujfwnq8NgxeOsUsrGuK
TNltFhELjPhk9nf6N/xfOobBX8SU7OKC2ev6CkI6EpDSgZqySlqjZY80CI0WEivLap86JAgkdb3F
TF2tP/VGpD+jBtNLdQr1PHDz7KAZU4oGRfJioFg/0ZNOmKH/zYe4VEQ55UBQRTIN9+rf5tcGRE00
OIE4P2xMnrtuYd3unDh4vqnUg7+tBhwelx1qCaL0qosTjLhv3Tg3N1SS8gvt3Sh1g3MuN31rEk9D
I4a2ZIAnivAWifvE4DqAQo73pqxLBLJXkfD2gN6Uoe0MjiPLYiFjfd5+v2oKNdd+4JkT2HMTWAKB
DwOviheae2KfrCYFG+QENq/DvAKYE311U8DDXDD+qYW5QsjcEZ1YRH8lX0TIlWqzKTtDl+VMUYq1
TehLKuBjnD7jfkv6h+R1uBFidWOzAOLLhAHXhiNZVCLztpR/uxkUQvOQbGMBMcf6qLTG0k7NeWXm
L5CN7ptuCCFGoovRb9f6XWLHjTXmzE0UKGA0NzFfJaYZk6UbYslNDvV1BFwGuF5Ch1T9DMGabsAG
JSUyuzyAKFrAEzMeZouc0HCTiIxa7OlK+CsvD/0rndKjSMsgUN1n9aONwm1EpGuBzRWEBuNy/FBA
s/ME+d1slgswj/qX0pr5QF84MT81Qv5t8RDDnc7sNlxwp6JDeBUxgDJUh/enthzjvR6CIcDKOubm
BKw+mIBwRzfQfF7KImjFLLP1liH5f9RHey4bUSjrcVJwZDNpR+2b6ilD1KvwY47ZTzyf5rUcYLqs
ps75KSD3QEvCMoxNG+T0WuZ+g3Fw+s0Mk5CEkmLlD1P4CTx1Z55+H9h8+VoYzFYZrB50NW2w3CxJ
FJ+RRgIxhxGmhOaY/0NYuR51ZU5uy4/E6zq+u2YkLa8wl1ZOIr8sIzynB+zVx1jQcYVzNeyedSOG
b6CpTF08+kT6PDj3t1qZ7TI5VdnLB93cMHC+ORvs0rn0+HyWJM8SVyic0oT8gpRqjkumilia/7sg
rapeqOAqYA0I72oC868lRbAPosIB6Yub123V8EdRvA+scWbc+QxZm78ZyF9cVvOkj+J7EFe1zac1
O1U6XXJlwmERW8EldJnQsgB+Xz8FGLzmMtqy20zF9BEeRQ1KaiNe4wAZcmdwTkN1N/jUbGJhuerN
B7Z8teqhcUxNX6r1RbD6ZJHlND1eXebrll1UdkAPSuYL4nhfgwzLJJAk6J0wfahESwk+Ym/qDKSC
hiiTpzcAgMNmPL9L/MZeigHm5UtH96oidp5KozJb/gvCQpcG9SJ91171bXAFT4IgbnPYrJr4Tzsk
U1F8B5T0C3Blsyrh9Sm2/ROPlQive2jC+fIOZtMtUc4zhFyetEN6cjf4z4Ij7EWVkJ7hCNa/DcEe
XkCexuMIKrW/wrHJBytb141ga+hU63hy8gUomsDlFTsOxgpmBs9+fPlnRwFPLhOko30+BkbE4cw6
dBbVYvou9vdEcg/0jBS6PyPzY97UBQKYLXdp1EwEYXV5/NnXmbBu6ltreY5kyx6dawrTUL0eoNWb
1oh8BMuDaCp6vmZ7v1rS+6EUaRdLJStixjkplNcc/A8g3zNS6VGunP3GsHWQ+wf/7X8ULrlEj9Zr
Y5ace4W5D+TrZUXxGlgeQ2PBuoAXo9U2yk42ZeryV/0xb8rK3CIj8CPuGdSfFsSYxjhAtjr1LZcR
VQh1YEbjKXMeRkJRClLIOyS+tuezhiZ/+EJUBgg58WrwfVGE8fgGy2FgYUyrN1i0Ftfyw+C72O1t
a9KJTKyxbohMRDp9Pv+D9V9jWRwDM9pmNiCu8Csjlniv1obaMcLZAdf4LzPXmic7txg2RMQt8DlQ
sDxPkH0GTeDtP2jfyoGX8m7zYpHvnCXwMLC/jxhgaGm7kEN2T7bqDoqANShBMHVuuJ/HwNvvGyya
jcN/8yjGno47gTSaHuN2zfNUH7IOm0V7xEe/JRcGa2uGHr7uXGTL0cVHYqcxWXF9rpfxTow/Oyma
BraOMdptglKqoH20ueBIf/5jr/SWzGUJTe/HpaNXWZnQlLVunliP5S90PHsgt3LPWWho41hiR+Rt
ZVSbOzzWs23uCaDINeBhYewjgshL/GfISEVt3WArDCRKdf8bzA6OoxHEIX/1dHbvcXVwlitwn6P5
pYARkI8WIirqs2y22naukl4V1ALxrX1ntIk4CmmLiHmsbJ6brOfxFyyM179xadtvu0u5LmAz6AcF
FNQLHmYdvSeX1wWtAm82B5hjPGV71NvCrYTWeYs+mf/qXNAXH8L3hZDPn0vbU0Rbwmt2pr6VjkDR
pWXcBmrePqZlgx2VFv+gk3dTVUgdfn9b25uo2aVemIk2kVOMUPCKaBts8OLTUoOBt65Bn4CwFE1D
WwpzABqkrg3DlazQaEEH+QsVFOxjZgfZXU8b8wvBK7ZrmoIBJsexUnK3zw4BgThf8jO/TSIxzp1Y
Ih+5+IMmIPjJfGoloRoVt/DD/k6aOzI2t8VK8v667GhPoj7t/eP5fI+kbVxVKbkKrCC/0c/EKjgg
Uh6t0okNgtWZFRuHskvC2zTEKRs/NRVop7b4CXpkkBz6qcs39LVeFG8lNz/CMyC/ZZ2sAiy4RpnC
KsIt8asGdRNfzGLoFn9A5hn7bk6mKZAj7zUwisqUUfnWPtLfi8WsMs7y/hCEioYWj5M6dDF2YV2S
31bi+a/EDLGS2UqF+nvMjuKXv9KHUWEAWe95tXUg5m17g0xJhqlhYVV5alq7ZOgMNPlox8A+2U8b
KZjFJQ==
`protect end_protected
